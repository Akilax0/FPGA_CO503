// SoC.v

// Generated using ACDS version 12.1 177 at 2022.03.30.07:47:41

`timescale 1 ps / 1 ps
module SoC (
		input  wire  reset_reset_n, // reset.reset_n
		input  wire  clk_clk        //   clk.clk
	);

	wire         cpu0_instruction_master_waitrequest;                                                                // cpu0_instruction_master_translator:av_waitrequest -> cpu0:i_waitrequest
	wire  [17:0] cpu0_instruction_master_address;                                                                    // cpu0:i_address -> cpu0_instruction_master_translator:av_address
	wire         cpu0_instruction_master_read;                                                                       // cpu0:i_read -> cpu0_instruction_master_translator:av_read
	wire  [31:0] cpu0_instruction_master_readdata;                                                                   // cpu0_instruction_master_translator:av_readdata -> cpu0:i_readdata
	wire         cpu0_instruction_master_readdatavalid;                                                              // cpu0_instruction_master_translator:av_readdatavalid -> cpu0:i_readdatavalid
	wire         cpu0_data_master_waitrequest;                                                                       // cpu0_data_master_translator:av_waitrequest -> cpu0:d_waitrequest
	wire  [31:0] cpu0_data_master_writedata;                                                                         // cpu0:d_writedata -> cpu0_data_master_translator:av_writedata
	wire  [17:0] cpu0_data_master_address;                                                                           // cpu0:d_address -> cpu0_data_master_translator:av_address
	wire         cpu0_data_master_write;                                                                             // cpu0:d_write -> cpu0_data_master_translator:av_write
	wire         cpu0_data_master_read;                                                                              // cpu0:d_read -> cpu0_data_master_translator:av_read
	wire  [31:0] cpu0_data_master_readdata;                                                                          // cpu0_data_master_translator:av_readdata -> cpu0:d_readdata
	wire         cpu0_data_master_debugaccess;                                                                       // cpu0:jtag_debug_module_debugaccess_to_roms -> cpu0_data_master_translator:av_debugaccess
	wire   [3:0] cpu0_data_master_byteenable;                                                                        // cpu0:d_byteenable -> cpu0_data_master_translator:av_byteenable
	wire         cpu1_data_master_waitrequest;                                                                       // cpu1_data_master_translator:av_waitrequest -> cpu1:d_waitrequest
	wire  [31:0] cpu1_data_master_writedata;                                                                         // cpu1:d_writedata -> cpu1_data_master_translator:av_writedata
	wire  [17:0] cpu1_data_master_address;                                                                           // cpu1:d_address -> cpu1_data_master_translator:av_address
	wire         cpu1_data_master_write;                                                                             // cpu1:d_write -> cpu1_data_master_translator:av_write
	wire         cpu1_data_master_read;                                                                              // cpu1:d_read -> cpu1_data_master_translator:av_read
	wire  [31:0] cpu1_data_master_readdata;                                                                          // cpu1_data_master_translator:av_readdata -> cpu1:d_readdata
	wire         cpu1_data_master_debugaccess;                                                                       // cpu1:jtag_debug_module_debugaccess_to_roms -> cpu1_data_master_translator:av_debugaccess
	wire   [3:0] cpu1_data_master_byteenable;                                                                        // cpu1:d_byteenable -> cpu1_data_master_translator:av_byteenable
	wire         cpu1_instruction_master_waitrequest;                                                                // cpu1_instruction_master_translator:av_waitrequest -> cpu1:i_waitrequest
	wire  [17:0] cpu1_instruction_master_address;                                                                    // cpu1:i_address -> cpu1_instruction_master_translator:av_address
	wire         cpu1_instruction_master_read;                                                                       // cpu1:i_read -> cpu1_instruction_master_translator:av_read
	wire  [31:0] cpu1_instruction_master_readdata;                                                                   // cpu1_instruction_master_translator:av_readdata -> cpu1:i_readdata
	wire         cpu1_instruction_master_readdatavalid;                                                              // cpu1_instruction_master_translator:av_readdatavalid -> cpu1:i_readdatavalid
	wire  [31:0] cpu0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                    // cpu0_jtag_debug_module_translator:av_writedata -> cpu0:jtag_debug_module_writedata
	wire   [8:0] cpu0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                      // cpu0_jtag_debug_module_translator:av_address -> cpu0:jtag_debug_module_address
	wire         cpu0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                   // cpu0_jtag_debug_module_translator:av_chipselect -> cpu0:jtag_debug_module_select
	wire         cpu0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                        // cpu0_jtag_debug_module_translator:av_write -> cpu0:jtag_debug_module_write
	wire  [31:0] cpu0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                     // cpu0:jtag_debug_module_readdata -> cpu0_jtag_debug_module_translator:av_readdata
	wire         cpu0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                // cpu0_jtag_debug_module_translator:av_begintransfer -> cpu0:jtag_debug_module_begintransfer
	wire         cpu0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                  // cpu0_jtag_debug_module_translator:av_debugaccess -> cpu0:jtag_debug_module_debugaccess
	wire   [3:0] cpu0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                   // cpu0_jtag_debug_module_translator:av_byteenable -> cpu0:jtag_debug_module_byteenable
	wire  [31:0] ins_mem0_s1_translator_avalon_anti_slave_0_writedata;                                               // ins_mem0_s1_translator:av_writedata -> ins_mem0:writedata
	wire  [13:0] ins_mem0_s1_translator_avalon_anti_slave_0_address;                                                 // ins_mem0_s1_translator:av_address -> ins_mem0:address
	wire         ins_mem0_s1_translator_avalon_anti_slave_0_chipselect;                                              // ins_mem0_s1_translator:av_chipselect -> ins_mem0:chipselect
	wire         ins_mem0_s1_translator_avalon_anti_slave_0_clken;                                                   // ins_mem0_s1_translator:av_clken -> ins_mem0:clken
	wire         ins_mem0_s1_translator_avalon_anti_slave_0_write;                                                   // ins_mem0_s1_translator:av_write -> ins_mem0:write
	wire  [31:0] ins_mem0_s1_translator_avalon_anti_slave_0_readdata;                                                // ins_mem0:readdata -> ins_mem0_s1_translator:av_readdata
	wire   [3:0] ins_mem0_s1_translator_avalon_anti_slave_0_byteenable;                                              // ins_mem0_s1_translator:av_byteenable -> ins_mem0:byteenable
	wire  [31:0] data_mem0_s1_translator_avalon_anti_slave_0_writedata;                                              // data_mem0_s1_translator:av_writedata -> data_mem0:writedata
	wire  [12:0] data_mem0_s1_translator_avalon_anti_slave_0_address;                                                // data_mem0_s1_translator:av_address -> data_mem0:address
	wire         data_mem0_s1_translator_avalon_anti_slave_0_chipselect;                                             // data_mem0_s1_translator:av_chipselect -> data_mem0:chipselect
	wire         data_mem0_s1_translator_avalon_anti_slave_0_clken;                                                  // data_mem0_s1_translator:av_clken -> data_mem0:clken
	wire         data_mem0_s1_translator_avalon_anti_slave_0_write;                                                  // data_mem0_s1_translator:av_write -> data_mem0:write
	wire  [31:0] data_mem0_s1_translator_avalon_anti_slave_0_readdata;                                               // data_mem0:readdata -> data_mem0_s1_translator:av_readdata
	wire   [3:0] data_mem0_s1_translator_avalon_anti_slave_0_byteenable;                                             // data_mem0_s1_translator:av_byteenable -> data_mem0:byteenable
	wire         fifo_0_in_translator_avalon_anti_slave_0_waitrequest;                                               // fifo_0:avalonmm_write_slave_waitrequest -> fifo_0_in_translator:av_waitrequest
	wire  [31:0] fifo_0_in_translator_avalon_anti_slave_0_writedata;                                                 // fifo_0_in_translator:av_writedata -> fifo_0:avalonmm_write_slave_writedata
	wire         fifo_0_in_translator_avalon_anti_slave_0_write;                                                     // fifo_0_in_translator:av_write -> fifo_0:avalonmm_write_slave_write
	wire  [31:0] fifo_0_in_csr_translator_avalon_anti_slave_0_writedata;                                             // fifo_0_in_csr_translator:av_writedata -> fifo_0:wrclk_control_slave_writedata
	wire   [2:0] fifo_0_in_csr_translator_avalon_anti_slave_0_address;                                               // fifo_0_in_csr_translator:av_address -> fifo_0:wrclk_control_slave_address
	wire         fifo_0_in_csr_translator_avalon_anti_slave_0_write;                                                 // fifo_0_in_csr_translator:av_write -> fifo_0:wrclk_control_slave_write
	wire         fifo_0_in_csr_translator_avalon_anti_slave_0_read;                                                  // fifo_0_in_csr_translator:av_read -> fifo_0:wrclk_control_slave_read
	wire  [31:0] fifo_0_in_csr_translator_avalon_anti_slave_0_readdata;                                              // fifo_0:wrclk_control_slave_readdata -> fifo_0_in_csr_translator:av_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                  // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                    // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire   [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                         // sysid_control_slave_translator:av_address -> sysid:address
	wire  [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                        // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire  [31:0] cpu1_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                    // cpu1_jtag_debug_module_translator:av_writedata -> cpu1:jtag_debug_module_writedata
	wire   [8:0] cpu1_jtag_debug_module_translator_avalon_anti_slave_0_address;                                      // cpu1_jtag_debug_module_translator:av_address -> cpu1:jtag_debug_module_address
	wire         cpu1_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                   // cpu1_jtag_debug_module_translator:av_chipselect -> cpu1:jtag_debug_module_select
	wire         cpu1_jtag_debug_module_translator_avalon_anti_slave_0_write;                                        // cpu1_jtag_debug_module_translator:av_write -> cpu1:jtag_debug_module_write
	wire  [31:0] cpu1_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                     // cpu1:jtag_debug_module_readdata -> cpu1_jtag_debug_module_translator:av_readdata
	wire         cpu1_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                // cpu1_jtag_debug_module_translator:av_begintransfer -> cpu1:jtag_debug_module_begintransfer
	wire         cpu1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                  // cpu1_jtag_debug_module_translator:av_debugaccess -> cpu1:jtag_debug_module_debugaccess
	wire   [3:0] cpu1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                   // cpu1_jtag_debug_module_translator:av_byteenable -> cpu1:jtag_debug_module_byteenable
	wire  [31:0] ins_mem1_s1_translator_avalon_anti_slave_0_writedata;                                               // ins_mem1_s1_translator:av_writedata -> ins_mem1:writedata
	wire  [13:0] ins_mem1_s1_translator_avalon_anti_slave_0_address;                                                 // ins_mem1_s1_translator:av_address -> ins_mem1:address
	wire         ins_mem1_s1_translator_avalon_anti_slave_0_chipselect;                                              // ins_mem1_s1_translator:av_chipselect -> ins_mem1:chipselect
	wire         ins_mem1_s1_translator_avalon_anti_slave_0_clken;                                                   // ins_mem1_s1_translator:av_clken -> ins_mem1:clken
	wire         ins_mem1_s1_translator_avalon_anti_slave_0_write;                                                   // ins_mem1_s1_translator:av_write -> ins_mem1:write
	wire  [31:0] ins_mem1_s1_translator_avalon_anti_slave_0_readdata;                                                // ins_mem1:readdata -> ins_mem1_s1_translator:av_readdata
	wire   [3:0] ins_mem1_s1_translator_avalon_anti_slave_0_byteenable;                                              // ins_mem1_s1_translator:av_byteenable -> ins_mem1:byteenable
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_1:av_waitrequest -> jtag_uart_1_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_1_avalon_jtag_slave_translator:av_writedata -> jtag_uart_1:av_writedata
	wire   [0:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_1_avalon_jtag_slave_translator:av_address -> jtag_uart_1:av_address
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_1_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_1:av_chipselect
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_1_avalon_jtag_slave_translator:av_write -> jtag_uart_1:av_write_n
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_1_avalon_jtag_slave_translator:av_read -> jtag_uart_1:av_read_n
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_1:av_readdata -> jtag_uart_1_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_1_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_1_s1_translator:av_writedata -> timer_1:writedata
	wire   [2:0] timer_1_s1_translator_avalon_anti_slave_0_address;                                                  // timer_1_s1_translator:av_address -> timer_1:address
	wire         timer_1_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	wire         timer_1_s1_translator_avalon_anti_slave_0_write;                                                    // timer_1_s1_translator:av_write -> timer_1:write_n
	wire  [15:0] timer_1_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_1:readdata -> timer_1_s1_translator:av_readdata
	wire         fifo_0_out_translator_avalon_anti_slave_0_waitrequest;                                              // fifo_0:avalonmm_read_slave_waitrequest -> fifo_0_out_translator:av_waitrequest
	wire         fifo_0_out_translator_avalon_anti_slave_0_read;                                                     // fifo_0_out_translator:av_read -> fifo_0:avalonmm_read_slave_read
	wire  [31:0] fifo_0_out_translator_avalon_anti_slave_0_readdata;                                                 // fifo_0:avalonmm_read_slave_readdata -> fifo_0_out_translator:av_readdata
	wire  [31:0] data_mem1_s1_translator_avalon_anti_slave_0_writedata;                                              // data_mem1_s1_translator:av_writedata -> data_mem1:writedata
	wire  [12:0] data_mem1_s1_translator_avalon_anti_slave_0_address;                                                // data_mem1_s1_translator:av_address -> data_mem1:address
	wire         data_mem1_s1_translator_avalon_anti_slave_0_chipselect;                                             // data_mem1_s1_translator:av_chipselect -> data_mem1:chipselect
	wire         data_mem1_s1_translator_avalon_anti_slave_0_clken;                                                  // data_mem1_s1_translator:av_clken -> data_mem1:clken
	wire         data_mem1_s1_translator_avalon_anti_slave_0_write;                                                  // data_mem1_s1_translator:av_write -> data_mem1:write
	wire  [31:0] data_mem1_s1_translator_avalon_anti_slave_0_readdata;                                               // data_mem1:readdata -> data_mem1_s1_translator:av_readdata
	wire   [3:0] data_mem1_s1_translator_avalon_anti_slave_0_byteenable;                                             // data_mem1_s1_translator:av_byteenable -> data_mem1:byteenable
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_waitrequest;                           // cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu0_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu0_instruction_master_translator_avalon_universal_master_0_burstcount;                            // cpu0_instruction_master_translator:uav_burstcount -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu0_instruction_master_translator_avalon_universal_master_0_writedata;                             // cpu0_instruction_master_translator:uav_writedata -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu0_instruction_master_translator_avalon_universal_master_0_address;                               // cpu0_instruction_master_translator:uav_address -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_lock;                                  // cpu0_instruction_master_translator:uav_lock -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_write;                                 // cpu0_instruction_master_translator:uav_write -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_read;                                  // cpu0_instruction_master_translator:uav_read -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu0_instruction_master_translator_avalon_universal_master_0_readdata;                              // cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu0_instruction_master_translator:uav_readdata
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_debugaccess;                           // cpu0_instruction_master_translator:uav_debugaccess -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu0_instruction_master_translator_avalon_universal_master_0_byteenable;                            // cpu0_instruction_master_translator:uav_byteenable -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                         // cpu0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu0_instruction_master_translator:uav_readdatavalid
	wire         cpu0_data_master_translator_avalon_universal_master_0_waitrequest;                                  // cpu0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu0_data_master_translator:uav_waitrequest
	wire   [2:0] cpu0_data_master_translator_avalon_universal_master_0_burstcount;                                   // cpu0_data_master_translator:uav_burstcount -> cpu0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu0_data_master_translator_avalon_universal_master_0_writedata;                                    // cpu0_data_master_translator:uav_writedata -> cpu0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu0_data_master_translator_avalon_universal_master_0_address;                                      // cpu0_data_master_translator:uav_address -> cpu0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu0_data_master_translator_avalon_universal_master_0_lock;                                         // cpu0_data_master_translator:uav_lock -> cpu0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu0_data_master_translator_avalon_universal_master_0_write;                                        // cpu0_data_master_translator:uav_write -> cpu0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu0_data_master_translator_avalon_universal_master_0_read;                                         // cpu0_data_master_translator:uav_read -> cpu0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu0_data_master_translator_avalon_universal_master_0_readdata;                                     // cpu0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu0_data_master_translator:uav_readdata
	wire         cpu0_data_master_translator_avalon_universal_master_0_debugaccess;                                  // cpu0_data_master_translator:uav_debugaccess -> cpu0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu0_data_master_translator_avalon_universal_master_0_byteenable;                                   // cpu0_data_master_translator:uav_byteenable -> cpu0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu0_data_master_translator_avalon_universal_master_0_readdatavalid;                                // cpu0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu0_data_master_translator:uav_readdatavalid
	wire         cpu1_data_master_translator_avalon_universal_master_0_waitrequest;                                  // cpu1_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu1_data_master_translator:uav_waitrequest
	wire   [2:0] cpu1_data_master_translator_avalon_universal_master_0_burstcount;                                   // cpu1_data_master_translator:uav_burstcount -> cpu1_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu1_data_master_translator_avalon_universal_master_0_writedata;                                    // cpu1_data_master_translator:uav_writedata -> cpu1_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu1_data_master_translator_avalon_universal_master_0_address;                                      // cpu1_data_master_translator:uav_address -> cpu1_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu1_data_master_translator_avalon_universal_master_0_lock;                                         // cpu1_data_master_translator:uav_lock -> cpu1_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu1_data_master_translator_avalon_universal_master_0_write;                                        // cpu1_data_master_translator:uav_write -> cpu1_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu1_data_master_translator_avalon_universal_master_0_read;                                         // cpu1_data_master_translator:uav_read -> cpu1_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu1_data_master_translator_avalon_universal_master_0_readdata;                                     // cpu1_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu1_data_master_translator:uav_readdata
	wire         cpu1_data_master_translator_avalon_universal_master_0_debugaccess;                                  // cpu1_data_master_translator:uav_debugaccess -> cpu1_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu1_data_master_translator_avalon_universal_master_0_byteenable;                                   // cpu1_data_master_translator:uav_byteenable -> cpu1_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu1_data_master_translator_avalon_universal_master_0_readdatavalid;                                // cpu1_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu1_data_master_translator:uav_readdatavalid
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_waitrequest;                           // cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu1_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu1_instruction_master_translator_avalon_universal_master_0_burstcount;                            // cpu1_instruction_master_translator:uav_burstcount -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu1_instruction_master_translator_avalon_universal_master_0_writedata;                             // cpu1_instruction_master_translator:uav_writedata -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu1_instruction_master_translator_avalon_universal_master_0_address;                               // cpu1_instruction_master_translator:uav_address -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_lock;                                  // cpu1_instruction_master_translator:uav_lock -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_write;                                 // cpu1_instruction_master_translator:uav_write -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_read;                                  // cpu1_instruction_master_translator:uav_read -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu1_instruction_master_translator_avalon_universal_master_0_readdata;                              // cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu1_instruction_master_translator:uav_readdata
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_debugaccess;                           // cpu1_instruction_master_translator:uav_debugaccess -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu1_instruction_master_translator_avalon_universal_master_0_byteenable;                            // cpu1_instruction_master_translator:uav_byteenable -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_readdatavalid;                         // cpu1_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu1_instruction_master_translator:uav_readdatavalid
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // cpu0_jtag_debug_module_translator:uav_waitrequest -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                      // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu0_jtag_debug_module_translator:uav_writedata
	wire  [17:0] cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                        // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu0_jtag_debug_module_translator:uav_address
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                          // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu0_jtag_debug_module_translator:uav_write
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                           // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu0_jtag_debug_module_translator:uav_lock
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                           // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu0_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                       // cpu0_jtag_debug_module_translator:uav_readdata -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // cpu0_jtag_debug_module_translator:uav_readdatavalid -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu0_jtag_debug_module_translator:uav_byteenable
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                    // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // ins_mem0_s1_translator:uav_waitrequest -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ins_mem0_s1_translator:uav_burstcount
	wire  [31:0] ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ins_mem0_s1_translator:uav_writedata
	wire  [17:0] ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_address -> ins_mem0_s1_translator:uav_address
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_write -> ins_mem0_s1_translator:uav_write
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ins_mem0_s1_translator:uav_lock
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_read -> ins_mem0_s1_translator:uav_read
	wire  [31:0] ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // ins_mem0_s1_translator:uav_readdata -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // ins_mem0_s1_translator:uav_readdatavalid -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ins_mem0_s1_translator:uav_debugaccess
	wire   [3:0] ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // ins_mem0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ins_mem0_s1_translator:uav_byteenable
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ins_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // data_mem0_s1_translator:uav_waitrequest -> data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> data_mem0_s1_translator:uav_burstcount
	wire  [31:0] data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> data_mem0_s1_translator:uav_writedata
	wire  [17:0] data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_address -> data_mem0_s1_translator:uav_address
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_write -> data_mem0_s1_translator:uav_write
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> data_mem0_s1_translator:uav_lock
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_read -> data_mem0_s1_translator:uav_read
	wire  [31:0] data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // data_mem0_s1_translator:uav_readdata -> data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // data_mem0_s1_translator:uav_readdatavalid -> data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> data_mem0_s1_translator:uav_debugaccess
	wire   [3:0] data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // data_mem0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> data_mem0_s1_translator:uav_byteenable
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // data_mem0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // data_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> data_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // data_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> data_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // data_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> data_mem0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // fifo_0_in_translator:uav_waitrequest -> fifo_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_in_translator:uav_burstcount
	wire  [31:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_in_translator:uav_writedata
	wire  [17:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_in_translator:uav_address
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_in_translator:uav_write
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_in_translator:uav_lock
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_in_translator:uav_read
	wire  [31:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // fifo_0_in_translator:uav_readdata -> fifo_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // fifo_0_in_translator:uav_readdatavalid -> fifo_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_in_translator:uav_debugaccess
	wire   [3:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_in_translator:uav_byteenable
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // fifo_0_in_csr_translator:uav_waitrequest -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_in_csr_translator:uav_burstcount
	wire  [31:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_in_csr_translator:uav_writedata
	wire  [17:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_in_csr_translator:uav_address
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_in_csr_translator:uav_write
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_in_csr_translator:uav_lock
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_in_csr_translator:uav_read
	wire  [31:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // fifo_0_in_csr_translator:uav_readdata -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // fifo_0_in_csr_translator:uav_readdatavalid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_in_csr_translator:uav_debugaccess
	wire   [3:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_in_csr_translator:uav_byteenable
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [17:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [17:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire  [17:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // cpu1_jtag_debug_module_translator:uav_waitrequest -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu1_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                      // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu1_jtag_debug_module_translator:uav_writedata
	wire  [17:0] cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                        // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu1_jtag_debug_module_translator:uav_address
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                          // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu1_jtag_debug_module_translator:uav_write
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                           // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu1_jtag_debug_module_translator:uav_lock
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                           // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu1_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                       // cpu1_jtag_debug_module_translator:uav_readdata -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // cpu1_jtag_debug_module_translator:uav_readdatavalid -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu1_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu1_jtag_debug_module_translator:uav_byteenable
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                    // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // ins_mem1_s1_translator:uav_waitrequest -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ins_mem1_s1_translator:uav_burstcount
	wire  [31:0] ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ins_mem1_s1_translator:uav_writedata
	wire  [17:0] ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_address -> ins_mem1_s1_translator:uav_address
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_write -> ins_mem1_s1_translator:uav_write
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ins_mem1_s1_translator:uav_lock
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_read -> ins_mem1_s1_translator:uav_read
	wire  [31:0] ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // ins_mem1_s1_translator:uav_readdata -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // ins_mem1_s1_translator:uav_readdatavalid -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ins_mem1_s1_translator:uav_debugaccess
	wire   [3:0] ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // ins_mem1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ins_mem1_s1_translator:uav_byteenable
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ins_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_1_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_1_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_1_avalon_jtag_slave_translator:uav_writedata
	wire  [17:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_1_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_1_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_1_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_1_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_1_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_1_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_1_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_1_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	wire  [17:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	wire   [3:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // fifo_0_out_translator:uav_waitrequest -> fifo_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // fifo_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_out_translator:uav_burstcount
	wire  [31:0] fifo_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // fifo_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_out_translator:uav_writedata
	wire  [17:0] fifo_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // fifo_0_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_out_translator:uav_address
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // fifo_0_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_out_translator:uav_write
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // fifo_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_out_translator:uav_lock
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // fifo_0_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_out_translator:uav_read
	wire  [31:0] fifo_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // fifo_0_out_translator:uav_readdata -> fifo_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // fifo_0_out_translator:uav_readdatavalid -> fifo_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // fifo_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_out_translator:uav_debugaccess
	wire   [3:0] fifo_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // fifo_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_out_translator:uav_byteenable
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // fifo_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // fifo_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // fifo_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // fifo_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // fifo_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // fifo_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] fifo_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // fifo_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // fifo_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // data_mem1_s1_translator:uav_waitrequest -> data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> data_mem1_s1_translator:uav_burstcount
	wire  [31:0] data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> data_mem1_s1_translator:uav_writedata
	wire  [17:0] data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_address -> data_mem1_s1_translator:uav_address
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_write -> data_mem1_s1_translator:uav_write
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> data_mem1_s1_translator:uav_lock
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_read -> data_mem1_s1_translator:uav_read
	wire  [31:0] data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // data_mem1_s1_translator:uav_readdata -> data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // data_mem1_s1_translator:uav_readdatavalid -> data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> data_mem1_s1_translator:uav_debugaccess
	wire   [3:0] data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // data_mem1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> data_mem1_s1_translator:uav_byteenable
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // data_mem1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // data_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> data_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // data_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> data_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // data_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> data_mem1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // cpu0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                        // cpu0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // cpu0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [92:0] cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                         // cpu0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router:sink_ready -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // cpu0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         cpu0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                               // cpu0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         cpu0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // cpu0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [92:0] cpu0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                // cpu0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         cpu0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_001:sink_ready -> cpu0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // cpu1_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire         cpu1_data_master_translator_avalon_universal_master_0_agent_cp_valid;                               // cpu1_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire         cpu1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // cpu1_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [92:0] cpu1_data_master_translator_avalon_universal_master_0_agent_cp_data;                                // cpu1_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire         cpu1_data_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_002:sink_ready -> cpu1_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // cpu1_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                        // cpu1_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // cpu1_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [92:0] cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                         // cpu1_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire         cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_003:sink_ready -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                          // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [92:0] cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                           // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router:sink_ready -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [92:0] ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // ins_mem0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_001:sink_ready -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // data_mem0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // data_mem0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // data_mem0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [92:0] data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // data_mem0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_002:sink_ready -> data_mem0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // fifo_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // fifo_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // fifo_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [92:0] fifo_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // fifo_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_003:sink_ready -> fifo_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [92:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_004:sink_ready -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [92:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [92:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_006:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [92:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_007:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                          // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [92:0] cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                           // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_008:sink_ready -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [92:0] ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // ins_mem1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_009:sink_ready -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [92:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_010:sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [92:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_011:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // fifo_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // fifo_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // fifo_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [92:0] fifo_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // fifo_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         fifo_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_012:sink_ready -> fifo_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // data_mem1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // data_mem1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // data_mem1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [92:0] data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // data_mem1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_013:sink_ready -> data_mem1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                        // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                              // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                      // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [92:0] addr_router_src_data;                                                                               // addr_router:src_data -> limiter:cmd_sink_data
	wire  [13:0] addr_router_src_channel;                                                                            // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                              // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                        // limiter:rsp_src_endofpacket -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                              // limiter:rsp_src_valid -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                      // limiter:rsp_src_startofpacket -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [92:0] limiter_rsp_src_data;                                                                               // limiter:rsp_src_data -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [13:0] limiter_rsp_src_channel;                                                                            // limiter:rsp_src_channel -> cpu0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                              // cpu0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_003_src_endofpacket;                                                                    // addr_router_003:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_003_src_valid;                                                                          // addr_router_003:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_003_src_startofpacket;                                                                  // addr_router_003:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [92:0] addr_router_003_src_data;                                                                           // addr_router_003:src_data -> limiter_001:cmd_sink_data
	wire  [13:0] addr_router_003_src_channel;                                                                        // addr_router_003:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_003_src_ready;                                                                          // limiter_001:cmd_sink_ready -> addr_router_003:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                    // limiter_001:rsp_src_endofpacket -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                          // limiter_001:rsp_src_valid -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                  // limiter_001:rsp_src_startofpacket -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [92:0] limiter_001_rsp_src_data;                                                                           // limiter_001:rsp_src_data -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [13:0] limiter_001_rsp_src_channel;                                                                        // limiter_001:rsp_src_channel -> cpu1_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                          // cpu1_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         rst_controller_reset_out_reset;                                                                     // rst_controller:reset_out -> [cmd_xbar_mux_001:reset, id_router_001:reset, id_router_005:reset, id_router_006:reset, ins_mem0:reset, ins_mem0_s1_translator:reset, ins_mem0_s1_translator_avalon_universal_slave_0_agent:reset, ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cpu0_jtag_debug_module_reset_reset;                                                                 // cpu0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_003:reset_in2]
	wire         rst_controller_001_reset_out_reset;                                                                 // rst_controller_001:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_008:reset, cpu0:reset_n, cpu0_data_master_translator:reset, cpu0_data_master_translator_avalon_universal_master_0_agent:reset, cpu0_instruction_master_translator:reset, cpu0_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu0_jtag_debug_module_translator:reset, cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu1:reset_n, cpu1_data_master_translator:reset, cpu1_data_master_translator_avalon_universal_master_0_agent:reset, cpu1_instruction_master_translator:reset, cpu1_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu1_jtag_debug_module_translator:reset, cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, data_mem0:reset, data_mem0_s1_translator:reset, data_mem0_s1_translator_avalon_universal_slave_0_agent:reset, data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_002:reset, id_router_008:reset, irq_mapper:reset, irq_mapper_001:reset, limiter:reset, limiter_001:reset, rsp_xbar_demux:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_008:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, rsp_xbar_mux_003:reset]
	wire         rst_controller_002_reset_out_reset;                                                                 // rst_controller_002:reset_out -> [cmd_xbar_mux_007:reset, cmd_xbar_mux_009:reset, cmd_xbar_mux_013:reset, data_mem1:reset, data_mem1_s1_translator:reset, data_mem1_s1_translator_avalon_universal_slave_0_agent:reset, data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_007:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_013:reset, ins_mem1:reset, ins_mem1_s1_translator:reset, ins_mem1_s1_translator_avalon_universal_slave_0_agent:reset, ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, jtag_uart_1:rst_n, jtag_uart_1_avalon_jtag_slave_translator:reset, jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_013:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1:reset_n, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cpu1_jtag_debug_module_reset_reset;                                                                 // cpu1:jtag_debug_module_resetrequest -> [rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_003_reset_out_reset;                                                                 // rst_controller_003:reset_out -> [cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_012:reset, fifo_0:reset_n, fifo_0_in_csr_translator:reset, fifo_0_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_in_translator:reset, fifo_0_in_translator_avalon_universal_slave_0_agent:reset, fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_out_translator:reset, fifo_0_out_translator_avalon_universal_slave_0_agent:reset, fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_003:reset, id_router_004:reset, id_router_012:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_012:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                    // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                          // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                  // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_src0_data;                                                                           // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [13:0] cmd_xbar_demux_src0_channel;                                                                        // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                          // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                    // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                          // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                  // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_src1_data;                                                                           // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [13:0] cmd_xbar_demux_src1_channel;                                                                        // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                          // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                    // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                          // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                  // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_src2_data;                                                                           // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [13:0] cmd_xbar_demux_src2_channel;                                                                        // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                          // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                    // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                          // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                  // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_src3_data;                                                                           // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire  [13:0] cmd_xbar_demux_src3_channel;                                                                        // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                          // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_src4_endofpacket;                                                                    // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                          // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                  // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_src4_data;                                                                           // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire  [13:0] cmd_xbar_demux_src4_channel;                                                                        // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire         cmd_xbar_demux_src4_ready;                                                                          // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                      // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                              // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src0_data;                                                                       // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [13:0] cmd_xbar_demux_001_src0_channel;                                                                    // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                      // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                      // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                              // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src1_data;                                                                       // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [13:0] cmd_xbar_demux_001_src1_channel;                                                                    // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                      // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                      // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                              // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src2_data;                                                                       // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [13:0] cmd_xbar_demux_001_src2_channel;                                                                    // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                      // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                      // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                              // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src3_data;                                                                       // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire  [13:0] cmd_xbar_demux_001_src3_channel;                                                                    // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                      // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                      // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                              // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src4_data;                                                                       // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire  [13:0] cmd_xbar_demux_001_src4_channel;                                                                    // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire         cmd_xbar_demux_001_src4_ready;                                                                      // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                // cmd_xbar_demux_001:src5_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                      // cmd_xbar_demux_001:src5_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                              // cmd_xbar_demux_001:src5_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src5_data;                                                                       // cmd_xbar_demux_001:src5_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src5_channel;                                                                    // cmd_xbar_demux_001:src5_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                // cmd_xbar_demux_001:src6_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                      // cmd_xbar_demux_001:src6_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                              // cmd_xbar_demux_001:src6_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src6_data;                                                                       // cmd_xbar_demux_001:src6_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src6_channel;                                                                    // cmd_xbar_demux_001:src6_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                // cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                      // cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink0_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                              // cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src7_data;                                                                       // cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink0_data
	wire  [13:0] cmd_xbar_demux_001_src7_channel;                                                                    // cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink0_channel
	wire         cmd_xbar_demux_001_src7_ready;                                                                      // cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux_001:src7_ready
	wire         cmd_xbar_demux_002_src0_endofpacket;                                                                // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire         cmd_xbar_demux_002_src0_valid;                                                                      // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_007:sink1_valid
	wire         cmd_xbar_demux_002_src0_startofpacket;                                                              // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_002_src0_data;                                                                       // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_007:sink1_data
	wire  [13:0] cmd_xbar_demux_002_src0_channel;                                                                    // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_007:sink1_channel
	wire         cmd_xbar_demux_002_src0_ready;                                                                      // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire         cmd_xbar_demux_002_src1_endofpacket;                                                                // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire         cmd_xbar_demux_002_src1_valid;                                                                      // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_008:sink0_valid
	wire         cmd_xbar_demux_002_src1_startofpacket;                                                              // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_002_src1_data;                                                                       // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_008:sink0_data
	wire  [13:0] cmd_xbar_demux_002_src1_channel;                                                                    // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_008:sink0_channel
	wire         cmd_xbar_demux_002_src1_ready;                                                                      // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux_002:src1_ready
	wire         cmd_xbar_demux_002_src2_endofpacket;                                                                // cmd_xbar_demux_002:src2_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire         cmd_xbar_demux_002_src2_valid;                                                                      // cmd_xbar_demux_002:src2_valid -> cmd_xbar_mux_009:sink0_valid
	wire         cmd_xbar_demux_002_src2_startofpacket;                                                              // cmd_xbar_demux_002:src2_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_002_src2_data;                                                                       // cmd_xbar_demux_002:src2_data -> cmd_xbar_mux_009:sink0_data
	wire  [13:0] cmd_xbar_demux_002_src2_channel;                                                                    // cmd_xbar_demux_002:src2_channel -> cmd_xbar_mux_009:sink0_channel
	wire         cmd_xbar_demux_002_src2_ready;                                                                      // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux_002:src2_ready
	wire         cmd_xbar_demux_002_src3_endofpacket;                                                                // cmd_xbar_demux_002:src3_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src3_valid;                                                                      // cmd_xbar_demux_002:src3_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src3_startofpacket;                                                              // cmd_xbar_demux_002:src3_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_002_src3_data;                                                                       // cmd_xbar_demux_002:src3_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_002_src3_channel;                                                                    // cmd_xbar_demux_002:src3_channel -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src4_endofpacket;                                                                // cmd_xbar_demux_002:src4_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src4_valid;                                                                      // cmd_xbar_demux_002:src4_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src4_startofpacket;                                                              // cmd_xbar_demux_002:src4_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_002_src4_data;                                                                       // cmd_xbar_demux_002:src4_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_002_src4_channel;                                                                    // cmd_xbar_demux_002:src4_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src5_endofpacket;                                                                // cmd_xbar_demux_002:src5_endofpacket -> cmd_xbar_mux_012:sink0_endofpacket
	wire         cmd_xbar_demux_002_src5_valid;                                                                      // cmd_xbar_demux_002:src5_valid -> cmd_xbar_mux_012:sink0_valid
	wire         cmd_xbar_demux_002_src5_startofpacket;                                                              // cmd_xbar_demux_002:src5_startofpacket -> cmd_xbar_mux_012:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_002_src5_data;                                                                       // cmd_xbar_demux_002:src5_data -> cmd_xbar_mux_012:sink0_data
	wire  [13:0] cmd_xbar_demux_002_src5_channel;                                                                    // cmd_xbar_demux_002:src5_channel -> cmd_xbar_mux_012:sink0_channel
	wire         cmd_xbar_demux_002_src5_ready;                                                                      // cmd_xbar_mux_012:sink0_ready -> cmd_xbar_demux_002:src5_ready
	wire         cmd_xbar_demux_002_src6_endofpacket;                                                                // cmd_xbar_demux_002:src6_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	wire         cmd_xbar_demux_002_src6_valid;                                                                      // cmd_xbar_demux_002:src6_valid -> cmd_xbar_mux_013:sink0_valid
	wire         cmd_xbar_demux_002_src6_startofpacket;                                                              // cmd_xbar_demux_002:src6_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_002_src6_data;                                                                       // cmd_xbar_demux_002:src6_data -> cmd_xbar_mux_013:sink0_data
	wire  [13:0] cmd_xbar_demux_002_src6_channel;                                                                    // cmd_xbar_demux_002:src6_channel -> cmd_xbar_mux_013:sink0_channel
	wire         cmd_xbar_demux_002_src6_ready;                                                                      // cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux_002:src6_ready
	wire         cmd_xbar_demux_003_src0_endofpacket;                                                                // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire         cmd_xbar_demux_003_src0_valid;                                                                      // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_008:sink1_valid
	wire         cmd_xbar_demux_003_src0_startofpacket;                                                              // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_003_src0_data;                                                                       // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_008:sink1_data
	wire  [13:0] cmd_xbar_demux_003_src0_channel;                                                                    // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_008:sink1_channel
	wire         cmd_xbar_demux_003_src0_ready;                                                                      // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_003:src0_ready
	wire         cmd_xbar_demux_003_src1_endofpacket;                                                                // cmd_xbar_demux_003:src1_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire         cmd_xbar_demux_003_src1_valid;                                                                      // cmd_xbar_demux_003:src1_valid -> cmd_xbar_mux_009:sink1_valid
	wire         cmd_xbar_demux_003_src1_startofpacket;                                                              // cmd_xbar_demux_003:src1_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_003_src1_data;                                                                       // cmd_xbar_demux_003:src1_data -> cmd_xbar_mux_009:sink1_data
	wire  [13:0] cmd_xbar_demux_003_src1_channel;                                                                    // cmd_xbar_demux_003:src1_channel -> cmd_xbar_mux_009:sink1_channel
	wire         cmd_xbar_demux_003_src1_ready;                                                                      // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_003:src1_ready
	wire         cmd_xbar_demux_003_src2_endofpacket;                                                                // cmd_xbar_demux_003:src2_endofpacket -> cmd_xbar_mux_012:sink1_endofpacket
	wire         cmd_xbar_demux_003_src2_valid;                                                                      // cmd_xbar_demux_003:src2_valid -> cmd_xbar_mux_012:sink1_valid
	wire         cmd_xbar_demux_003_src2_startofpacket;                                                              // cmd_xbar_demux_003:src2_startofpacket -> cmd_xbar_mux_012:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_003_src2_data;                                                                       // cmd_xbar_demux_003:src2_data -> cmd_xbar_mux_012:sink1_data
	wire  [13:0] cmd_xbar_demux_003_src2_channel;                                                                    // cmd_xbar_demux_003:src2_channel -> cmd_xbar_mux_012:sink1_channel
	wire         cmd_xbar_demux_003_src2_ready;                                                                      // cmd_xbar_mux_012:sink1_ready -> cmd_xbar_demux_003:src2_ready
	wire         cmd_xbar_demux_003_src3_endofpacket;                                                                // cmd_xbar_demux_003:src3_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	wire         cmd_xbar_demux_003_src3_valid;                                                                      // cmd_xbar_demux_003:src3_valid -> cmd_xbar_mux_013:sink1_valid
	wire         cmd_xbar_demux_003_src3_startofpacket;                                                              // cmd_xbar_demux_003:src3_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_003_src3_data;                                                                       // cmd_xbar_demux_003:src3_data -> cmd_xbar_mux_013:sink1_data
	wire  [13:0] cmd_xbar_demux_003_src3_channel;                                                                    // cmd_xbar_demux_003:src3_channel -> cmd_xbar_mux_013:sink1_channel
	wire         cmd_xbar_demux_003_src3_ready;                                                                      // cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_003:src3_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                    // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                          // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                  // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [92:0] rsp_xbar_demux_src0_data;                                                                           // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [13:0] rsp_xbar_demux_src0_channel;                                                                        // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                          // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                    // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                          // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                  // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [92:0] rsp_xbar_demux_src1_data;                                                                           // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [13:0] rsp_xbar_demux_src1_channel;                                                                        // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                          // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                      // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                              // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [92:0] rsp_xbar_demux_001_src0_data;                                                                       // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [13:0] rsp_xbar_demux_001_src0_channel;                                                                    // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                      // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                      // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                              // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [92:0] rsp_xbar_demux_001_src1_data;                                                                       // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [13:0] rsp_xbar_demux_001_src1_channel;                                                                    // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                      // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                      // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                              // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [92:0] rsp_xbar_demux_002_src0_data;                                                                       // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [13:0] rsp_xbar_demux_002_src0_channel;                                                                    // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                      // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                      // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                              // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [92:0] rsp_xbar_demux_002_src1_data;                                                                       // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [13:0] rsp_xbar_demux_002_src1_channel;                                                                    // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                      // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                      // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                              // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [92:0] rsp_xbar_demux_003_src0_data;                                                                       // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire  [13:0] rsp_xbar_demux_003_src0_channel;                                                                    // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                      // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                                // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                      // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                              // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [92:0] rsp_xbar_demux_003_src1_data;                                                                       // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire  [13:0] rsp_xbar_demux_003_src1_channel;                                                                    // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                      // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                      // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                              // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [92:0] rsp_xbar_demux_004_src0_data;                                                                       // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire  [13:0] rsp_xbar_demux_004_src0_channel;                                                                    // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                      // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_004_src1_endofpacket;                                                                // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src1_valid;                                                                      // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src1_startofpacket;                                                              // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [92:0] rsp_xbar_demux_004_src1_data;                                                                       // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire  [13:0] rsp_xbar_demux_004_src1_channel;                                                                    // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src1_ready;                                                                      // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                      // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                              // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [92:0] rsp_xbar_demux_005_src0_data;                                                                       // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [13:0] rsp_xbar_demux_005_src0_channel;                                                                    // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                      // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                      // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                              // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [92:0] rsp_xbar_demux_006_src0_data;                                                                       // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [13:0] rsp_xbar_demux_006_src0_channel;                                                                    // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                      // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                      // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                              // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [92:0] rsp_xbar_demux_007_src0_data;                                                                       // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [13:0] rsp_xbar_demux_007_src0_channel;                                                                    // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                      // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_007_src1_endofpacket;                                                                // rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire         rsp_xbar_demux_007_src1_valid;                                                                      // rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_002:sink0_valid
	wire         rsp_xbar_demux_007_src1_startofpacket;                                                              // rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [92:0] rsp_xbar_demux_007_src1_data;                                                                       // rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_002:sink0_data
	wire  [13:0] rsp_xbar_demux_007_src1_channel;                                                                    // rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_002:sink0_channel
	wire         rsp_xbar_demux_007_src1_ready;                                                                      // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_007:src1_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                      // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_002:sink1_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                              // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [92:0] rsp_xbar_demux_008_src0_data;                                                                       // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_002:sink1_data
	wire  [13:0] rsp_xbar_demux_008_src0_channel;                                                                    // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_002:sink1_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                      // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_008_src1_endofpacket;                                                                // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire         rsp_xbar_demux_008_src1_valid;                                                                      // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_003:sink0_valid
	wire         rsp_xbar_demux_008_src1_startofpacket;                                                              // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [92:0] rsp_xbar_demux_008_src1_data;                                                                       // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_003:sink0_data
	wire  [13:0] rsp_xbar_demux_008_src1_channel;                                                                    // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_003:sink0_channel
	wire         rsp_xbar_demux_008_src1_ready;                                                                      // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_008:src1_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                      // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_002:sink2_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                              // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [92:0] rsp_xbar_demux_009_src0_data;                                                                       // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_002:sink2_data
	wire  [13:0] rsp_xbar_demux_009_src0_channel;                                                                    // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_002:sink2_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                      // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_009_src1_endofpacket;                                                                // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire         rsp_xbar_demux_009_src1_valid;                                                                      // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_003:sink1_valid
	wire         rsp_xbar_demux_009_src1_startofpacket;                                                              // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [92:0] rsp_xbar_demux_009_src1_data;                                                                       // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_003:sink1_data
	wire  [13:0] rsp_xbar_demux_009_src1_channel;                                                                    // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_003:sink1_channel
	wire         rsp_xbar_demux_009_src1_ready;                                                                      // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_009:src1_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                      // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_002:sink3_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                              // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [92:0] rsp_xbar_demux_010_src0_data;                                                                       // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_002:sink3_data
	wire  [13:0] rsp_xbar_demux_010_src0_channel;                                                                    // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_002:sink3_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                      // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                                // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                      // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_002:sink4_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                              // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	wire  [92:0] rsp_xbar_demux_011_src0_data;                                                                       // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_002:sink4_data
	wire  [13:0] rsp_xbar_demux_011_src0_channel;                                                                    // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_002:sink4_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                      // rsp_xbar_mux_002:sink4_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                                // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_002:sink5_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                      // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_002:sink5_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                              // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_002:sink5_startofpacket
	wire  [92:0] rsp_xbar_demux_012_src0_data;                                                                       // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_002:sink5_data
	wire  [13:0] rsp_xbar_demux_012_src0_channel;                                                                    // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_002:sink5_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                      // rsp_xbar_mux_002:sink5_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_012_src1_endofpacket;                                                                // rsp_xbar_demux_012:src1_endofpacket -> rsp_xbar_mux_003:sink2_endofpacket
	wire         rsp_xbar_demux_012_src1_valid;                                                                      // rsp_xbar_demux_012:src1_valid -> rsp_xbar_mux_003:sink2_valid
	wire         rsp_xbar_demux_012_src1_startofpacket;                                                              // rsp_xbar_demux_012:src1_startofpacket -> rsp_xbar_mux_003:sink2_startofpacket
	wire  [92:0] rsp_xbar_demux_012_src1_data;                                                                       // rsp_xbar_demux_012:src1_data -> rsp_xbar_mux_003:sink2_data
	wire  [13:0] rsp_xbar_demux_012_src1_channel;                                                                    // rsp_xbar_demux_012:src1_channel -> rsp_xbar_mux_003:sink2_channel
	wire         rsp_xbar_demux_012_src1_ready;                                                                      // rsp_xbar_mux_003:sink2_ready -> rsp_xbar_demux_012:src1_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                                // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_002:sink6_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                      // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_002:sink6_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                              // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_002:sink6_startofpacket
	wire  [92:0] rsp_xbar_demux_013_src0_data;                                                                       // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_002:sink6_data
	wire  [13:0] rsp_xbar_demux_013_src0_channel;                                                                    // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_002:sink6_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                      // rsp_xbar_mux_002:sink6_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_013_src1_endofpacket;                                                                // rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_003:sink3_endofpacket
	wire         rsp_xbar_demux_013_src1_valid;                                                                      // rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_003:sink3_valid
	wire         rsp_xbar_demux_013_src1_startofpacket;                                                              // rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_003:sink3_startofpacket
	wire  [92:0] rsp_xbar_demux_013_src1_data;                                                                       // rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_003:sink3_data
	wire  [13:0] rsp_xbar_demux_013_src1_channel;                                                                    // rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_003:sink3_channel
	wire         rsp_xbar_demux_013_src1_ready;                                                                      // rsp_xbar_mux_003:sink3_ready -> rsp_xbar_demux_013:src1_ready
	wire         limiter_cmd_src_endofpacket;                                                                        // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                      // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [92:0] limiter_cmd_src_data;                                                                               // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [13:0] limiter_cmd_src_channel;                                                                            // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                              // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                       // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                             // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                     // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [92:0] rsp_xbar_mux_src_data;                                                                              // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [13:0] rsp_xbar_mux_src_channel;                                                                           // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                             // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                    // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                          // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                  // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [92:0] addr_router_001_src_data;                                                                           // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire  [13:0] addr_router_001_src_channel;                                                                        // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                          // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                   // rsp_xbar_mux_001:src_endofpacket -> cpu0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                         // rsp_xbar_mux_001:src_valid -> cpu0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                 // rsp_xbar_mux_001:src_startofpacket -> cpu0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [92:0] rsp_xbar_mux_001_src_data;                                                                          // rsp_xbar_mux_001:src_data -> cpu0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [13:0] rsp_xbar_mux_001_src_channel;                                                                       // rsp_xbar_mux_001:src_channel -> cpu0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                         // cpu0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         addr_router_002_src_endofpacket;                                                                    // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire         addr_router_002_src_valid;                                                                          // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire         addr_router_002_src_startofpacket;                                                                  // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [92:0] addr_router_002_src_data;                                                                           // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire  [13:0] addr_router_002_src_channel;                                                                        // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire         addr_router_002_src_ready;                                                                          // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire         rsp_xbar_mux_002_src_endofpacket;                                                                   // rsp_xbar_mux_002:src_endofpacket -> cpu1_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_002_src_valid;                                                                         // rsp_xbar_mux_002:src_valid -> cpu1_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_002_src_startofpacket;                                                                 // rsp_xbar_mux_002:src_startofpacket -> cpu1_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [92:0] rsp_xbar_mux_002_src_data;                                                                          // rsp_xbar_mux_002:src_data -> cpu1_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [13:0] rsp_xbar_mux_002_src_channel;                                                                       // rsp_xbar_mux_002:src_channel -> cpu1_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_002_src_ready;                                                                         // cpu1_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                    // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                  // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [92:0] limiter_001_cmd_src_data;                                                                           // limiter_001:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire  [13:0] limiter_001_cmd_src_channel;                                                                        // limiter_001:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                          // cmd_xbar_demux_003:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_003_src_endofpacket;                                                                   // rsp_xbar_mux_003:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_003_src_valid;                                                                         // rsp_xbar_mux_003:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_003_src_startofpacket;                                                                 // rsp_xbar_mux_003:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [92:0] rsp_xbar_mux_003_src_data;                                                                          // rsp_xbar_mux_003:src_data -> limiter_001:rsp_sink_data
	wire  [13:0] rsp_xbar_mux_003_src_channel;                                                                       // rsp_xbar_mux_003:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_003_src_ready;                                                                         // limiter_001:rsp_sink_ready -> rsp_xbar_mux_003:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                       // cmd_xbar_mux:src_endofpacket -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                             // cmd_xbar_mux:src_valid -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                     // cmd_xbar_mux:src_startofpacket -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_src_data;                                                                              // cmd_xbar_mux:src_data -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_src_channel;                                                                           // cmd_xbar_mux:src_channel -> cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                             // cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                          // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                        // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [92:0] id_router_src_data;                                                                                 // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [13:0] id_router_src_channel;                                                                              // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                   // cmd_xbar_mux_001:src_endofpacket -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                         // cmd_xbar_mux_001:src_valid -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                 // cmd_xbar_mux_001:src_startofpacket -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_001_src_data;                                                                          // cmd_xbar_mux_001:src_data -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_001_src_channel;                                                                       // cmd_xbar_mux_001:src_channel -> ins_mem0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                         // ins_mem0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                      // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                            // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                    // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [92:0] id_router_001_src_data;                                                                             // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [13:0] id_router_001_src_channel;                                                                          // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                   // cmd_xbar_mux_002:src_endofpacket -> data_mem0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                         // cmd_xbar_mux_002:src_valid -> data_mem0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                 // cmd_xbar_mux_002:src_startofpacket -> data_mem0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_002_src_data;                                                                          // cmd_xbar_mux_002:src_data -> data_mem0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_002_src_channel;                                                                       // cmd_xbar_mux_002:src_channel -> data_mem0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                         // data_mem0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                      // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                            // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                    // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [92:0] id_router_002_src_data;                                                                             // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [13:0] id_router_002_src_channel;                                                                          // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                   // cmd_xbar_mux_003:src_endofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                         // cmd_xbar_mux_003:src_valid -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                                 // cmd_xbar_mux_003:src_startofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_003_src_data;                                                                          // cmd_xbar_mux_003:src_data -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_003_src_channel;                                                                       // cmd_xbar_mux_003:src_channel -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                         // fifo_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire         id_router_003_src_endofpacket;                                                                      // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                            // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                    // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [92:0] id_router_003_src_data;                                                                             // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [13:0] id_router_003_src_channel;                                                                          // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_mux_004_src_endofpacket;                                                                   // cmd_xbar_mux_004:src_endofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_004_src_valid;                                                                         // cmd_xbar_mux_004:src_valid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_004_src_startofpacket;                                                                 // cmd_xbar_mux_004:src_startofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_004_src_data;                                                                          // cmd_xbar_mux_004:src_data -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_004_src_channel;                                                                       // cmd_xbar_mux_004:src_channel -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_004_src_ready;                                                                         // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire         id_router_004_src_endofpacket;                                                                      // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                            // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                    // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [92:0] id_router_004_src_data;                                                                             // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [13:0] id_router_004_src_channel;                                                                          // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                      // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                            // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                    // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [92:0] id_router_005_src_data;                                                                             // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [13:0] id_router_005_src_channel;                                                                          // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                            // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                      // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                            // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                    // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [92:0] id_router_006_src_data;                                                                             // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [13:0] id_router_006_src_channel;                                                                          // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                            // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_mux_007_src_endofpacket;                                                                   // cmd_xbar_mux_007:src_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_007_src_valid;                                                                         // cmd_xbar_mux_007:src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_007_src_startofpacket;                                                                 // cmd_xbar_mux_007:src_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_007_src_data;                                                                          // cmd_xbar_mux_007:src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_007_src_channel;                                                                       // cmd_xbar_mux_007:src_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_007_src_ready;                                                                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	wire         id_router_007_src_endofpacket;                                                                      // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                            // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                    // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [92:0] id_router_007_src_data;                                                                             // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [13:0] id_router_007_src_channel;                                                                          // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                            // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_mux_008_src_endofpacket;                                                                   // cmd_xbar_mux_008:src_endofpacket -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_008_src_valid;                                                                         // cmd_xbar_mux_008:src_valid -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_008_src_startofpacket;                                                                 // cmd_xbar_mux_008:src_startofpacket -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_008_src_data;                                                                          // cmd_xbar_mux_008:src_data -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_008_src_channel;                                                                       // cmd_xbar_mux_008:src_channel -> cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_008_src_ready;                                                                         // cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire         id_router_008_src_endofpacket;                                                                      // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                            // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                    // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [92:0] id_router_008_src_data;                                                                             // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [13:0] id_router_008_src_channel;                                                                          // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                            // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_mux_009_src_endofpacket;                                                                   // cmd_xbar_mux_009:src_endofpacket -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_009_src_valid;                                                                         // cmd_xbar_mux_009:src_valid -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_009_src_startofpacket;                                                                 // cmd_xbar_mux_009:src_startofpacket -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_009_src_data;                                                                          // cmd_xbar_mux_009:src_data -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_009_src_channel;                                                                       // cmd_xbar_mux_009:src_channel -> ins_mem1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_009_src_ready;                                                                         // ins_mem1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire         id_router_009_src_endofpacket;                                                                      // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                            // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                    // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [92:0] id_router_009_src_data;                                                                             // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [13:0] id_router_009_src_channel;                                                                          // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                            // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_demux_002_src3_ready;                                                                      // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src3_ready
	wire         id_router_010_src_endofpacket;                                                                      // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                            // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                    // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [92:0] id_router_010_src_data;                                                                             // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [13:0] id_router_010_src_channel;                                                                          // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                            // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_demux_002_src4_ready;                                                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src4_ready
	wire         id_router_011_src_endofpacket;                                                                      // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                            // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                    // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [92:0] id_router_011_src_data;                                                                             // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [13:0] id_router_011_src_channel;                                                                          // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                            // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_mux_012_src_endofpacket;                                                                   // cmd_xbar_mux_012:src_endofpacket -> fifo_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_012_src_valid;                                                                         // cmd_xbar_mux_012:src_valid -> fifo_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_012_src_startofpacket;                                                                 // cmd_xbar_mux_012:src_startofpacket -> fifo_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_012_src_data;                                                                          // cmd_xbar_mux_012:src_data -> fifo_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_012_src_channel;                                                                       // cmd_xbar_mux_012:src_channel -> fifo_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_012_src_ready;                                                                         // fifo_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_012:src_ready
	wire         id_router_012_src_endofpacket;                                                                      // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                            // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                    // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [92:0] id_router_012_src_data;                                                                             // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [13:0] id_router_012_src_channel;                                                                          // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                            // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_mux_013_src_endofpacket;                                                                   // cmd_xbar_mux_013:src_endofpacket -> data_mem1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_013_src_valid;                                                                         // cmd_xbar_mux_013:src_valid -> data_mem1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_013_src_startofpacket;                                                                 // cmd_xbar_mux_013:src_startofpacket -> data_mem1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_013_src_data;                                                                          // cmd_xbar_mux_013:src_data -> data_mem1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_013_src_channel;                                                                       // cmd_xbar_mux_013:src_channel -> data_mem1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_013_src_ready;                                                                         // data_mem1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	wire         id_router_013_src_endofpacket;                                                                      // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                            // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                    // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [92:0] id_router_013_src_data;                                                                             // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire  [13:0] id_router_013_src_channel;                                                                          // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                            // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire  [13:0] limiter_cmd_valid_data;                                                                             // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire  [13:0] limiter_001_cmd_valid_data;                                                                         // limiter_001:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                           // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                           // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu0_d_irq_irq;                                                                                     // irq_mapper:sender_irq -> cpu0:d_irq
	wire         irq_mapper_001_receiver0_irq;                                                                       // jtag_uart_1:av_irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                                                       // timer_1:irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] cpu1_d_irq_irq;                                                                                     // irq_mapper_001:sender_irq -> cpu1:d_irq
	wire         irq_mapper_receiver2_irq;                                                                           // fifo_0:wrclk_control_slave_irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver2_irq]

	SoC_ins_mem0 ins_mem0 (
		.clk        (clk_clk),                                               //   clk1.clk
		.address    (ins_mem0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ins_mem0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ins_mem0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ins_mem0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ins_mem0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ins_mem0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ins_mem0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                         // reset1.reset
	);

	SoC_cpu0 cpu0 (
		.clk                                   (clk_clk),                                                             //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                 //                   reset_n.reset_n
		.d_address                             (cpu0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu0_data_master_read),                                               //                          .read
		.d_readdata                            (cpu0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu0_data_master_write),                                              //                          .write
		.d_writedata                           (cpu0_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu0_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu0_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu0_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                     // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	SoC_timer_0 timer_0 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                              //   irq.irq
	);

	SoC_ins_mem1 ins_mem1 (
		.clk        (clk_clk),                                               //   clk1.clk
		.address    (ins_mem1_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ins_mem1_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ins_mem1_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ins_mem1_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ins_mem1_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ins_mem1_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ins_mem1_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset)                     // reset1.reset
	);

	SoC_cpu1 cpu1 (
		.clk                                   (clk_clk),                                                             //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                 //                   reset_n.reset_n
		.d_address                             (cpu1_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu1_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu1_data_master_read),                                               //                          .read
		.d_readdata                            (cpu1_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu1_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu1_data_master_write),                                              //                          .write
		.d_writedata                           (cpu1_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu1_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu1_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu1_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu1_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu1_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu1_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu1_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu1_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                     // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_1 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver0_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_1 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                  // reset.reset_n
		.address    (timer_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_001_receiver1_irq)                          //   irq.irq
	);

	SoC_sysid sysid (
		.clock    (clk_clk),                                                     //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	SoC_fifo_0 fifo_0 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_003_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (fifo_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver2_irq),                               //   in_irq.irq
		.avalonmm_read_slave_readdata     (fifo_0_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (fifo_0_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (fifo_0_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_data_mem0 data_mem0 (
		.clk        (clk_clk),                                                //   clk1.clk
		.address    (data_mem0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (data_mem0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (data_mem0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (data_mem0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (data_mem0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (data_mem0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (data_mem0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset)                      // reset1.reset
	);

	SoC_data_mem1 data_mem1 (
		.clk        (clk_clk),                                                //   clk1.clk
		.address    (data_mem1_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (data_mem1_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (data_mem1_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (data_mem1_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (data_mem1_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (data_mem1_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (data_mem1_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset)                      // reset1.reset
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu0_instruction_master_translator (
		.clk                   (clk_clk),                                                                    //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                         //                     reset.reset
		.uav_address           (cpu0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu0_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu0_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu0_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                       //               (terminated)
		.av_byteenable         (4'b1111),                                                                    //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                       //               (terminated)
		.av_begintransfer      (1'b0),                                                                       //               (terminated)
		.av_chipselect         (1'b0),                                                                       //               (terminated)
		.av_write              (1'b0),                                                                       //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                       //               (terminated)
		.av_lock               (1'b0),                                                                       //               (terminated)
		.av_debugaccess        (1'b0),                                                                       //               (terminated)
		.uav_clken             (),                                                                           //               (terminated)
		.av_clken              (1'b1)                                                                        //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu0_data_master_translator (
		.clk                   (clk_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                  //                     reset.reset
		.uav_address           (cpu0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu0_data_master_read),                                               //                          .read
		.av_readdata           (cpu0_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu0_data_master_write),                                              //                          .write
		.av_writedata          (cpu0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                //               (terminated)
		.av_begintransfer      (1'b0),                                                                //               (terminated)
		.av_chipselect         (1'b0),                                                                //               (terminated)
		.av_readdatavalid      (),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                //               (terminated)
		.uav_clken             (),                                                                    //               (terminated)
		.av_clken              (1'b1)                                                                 //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu1_data_master_translator (
		.clk                   (clk_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                  //                     reset.reset
		.uav_address           (cpu1_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu1_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu1_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu1_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu1_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu1_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu1_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu1_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu1_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu1_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu1_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu1_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu1_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu1_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu1_data_master_read),                                               //                          .read
		.av_readdata           (cpu1_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu1_data_master_write),                                              //                          .write
		.av_writedata          (cpu1_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu1_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                //               (terminated)
		.av_begintransfer      (1'b0),                                                                //               (terminated)
		.av_chipselect         (1'b0),                                                                //               (terminated)
		.av_readdatavalid      (),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                //               (terminated)
		.uav_clken             (),                                                                    //               (terminated)
		.av_clken              (1'b1)                                                                 //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu1_instruction_master_translator (
		.clk                   (clk_clk),                                                                    //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                         //                     reset.reset
		.uav_address           (cpu1_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu1_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu1_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu1_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu1_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu1_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu1_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu1_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu1_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu1_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu1_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu1_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu1_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu1_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu1_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu1_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                       //               (terminated)
		.av_byteenable         (4'b1111),                                                                    //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                       //               (terminated)
		.av_begintransfer      (1'b0),                                                                       //               (terminated)
		.av_chipselect         (1'b0),                                                                       //               (terminated)
		.av_write              (1'b0),                                                                       //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                       //               (terminated)
		.av_lock               (1'b0),                                                                       //               (terminated)
		.av_debugaccess        (1'b0),                                                                       //               (terminated)
		.uav_clken             (),                                                                           //               (terminated)
		.av_clken              (1'b1)                                                                        //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu0_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address           (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (14),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ins_mem0_s1_translator (
		.clk                   (clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ins_mem0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ins_mem0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ins_mem0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ins_mem0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ins_mem0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ins_mem0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ins_mem0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_mem0_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address           (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_mem0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (data_mem0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (data_mem0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (data_mem0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (data_mem0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (data_mem0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (data_mem0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                   //                    reset.reset
		.uav_address           (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (fifo_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (fifo_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                       //                    reset.reset
		.uav_address           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                             //                    reset.reset
		.uav_address           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_writedata          (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu1_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address           (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (14),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ins_mem1_s1_translator (
		.clk                   (clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                     //                    reset.reset
		.uav_address           (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ins_mem1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ins_mem1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ins_mem1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ins_mem1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ins_mem1_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ins_mem1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ins_mem1_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_1_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_1_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                    //                    reset.reset
		.uav_address           (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (fifo_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (fifo_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (fifo_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_mem1_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                      //                    reset.reset
		.uav_address           (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_mem1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (data_mem1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (data_mem1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (data_mem1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (data_mem1_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (data_mem1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (data_mem1_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (14),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                             //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.av_address       (cpu0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                               //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                             //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                         //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (14),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                      //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.av_address       (cpu0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                   //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                    //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                 //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                             //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                    //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (14),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu1_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                      //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.av_address       (cpu1_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu1_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu1_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu1_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu1_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu1_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu1_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu1_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu1_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu1_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu1_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_002_src_valid),                                                   //        rp.valid
		.rp_data          (rsp_xbar_mux_002_src_data),                                                    //          .data
		.rp_channel       (rsp_xbar_mux_002_src_channel),                                                 //          .channel
		.rp_startofpacket (rsp_xbar_mux_002_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_002_src_endofpacket),                                             //          .endofpacket
		.rp_ready         (rsp_xbar_mux_002_src_ready)                                                    //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (14),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu1_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                             //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.av_address       (cpu1_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu1_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu1_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu1_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu1_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu1_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu1_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu1_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu1_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu1_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu1_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                           //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                            //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                         //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                     //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                            //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                    //                .channel
		.rf_sink_ready           (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ins_mem0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ins_mem0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                     //                .channel
		.rf_sink_ready           (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_mem0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_mem0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                      //                .channel
		.rf_sink_ready           (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_mem0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_mem0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_mem0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                   //                .channel
		.rf_sink_ready           (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                             // clk_reset.reset
		.in_data           (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                       //                .channel
		.rf_sink_ready           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                 //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_007_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_007_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_007_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_007_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_007_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_007_src_channel),                                                             //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                                //                .channel
		.rf_sink_ready           (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ins_mem1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ins_mem1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                     //                .channel
		.rf_sink_ready           (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src3_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src3_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_002_src3_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src3_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src3_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src3_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src4_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src4_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src4_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src4_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src4_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src4_channel),                                                 //                .channel
		.rf_sink_ready           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_012_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_012_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_012_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_012_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_012_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_012_src_channel),                                                    //                .channel
		.rf_sink_ready           (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                              // clk_reset.reset
		.in_data           (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_mem1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_mem1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_013_src_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_mux_013_src_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_mux_013_src_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_mux_013_src_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_013_src_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_mux_013_src_channel),                                                      //                .channel
		.rf_sink_ready           (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_mem1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                // clk_reset.reset
		.in_data           (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_mem1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_mem1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	SoC_addr_router addr_router (
		.sink_ready         (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_src_valid),                                                               //          .valid
		.src_data           (addr_router_src_data),                                                                //          .data
		.src_channel        (addr_router_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                          //          .endofpacket
	);

	SoC_addr_router_001 addr_router_001 (
		.sink_ready         (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                    //          .valid
		.src_data           (addr_router_001_src_data),                                                     //          .data
		.src_channel        (addr_router_001_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                               //          .endofpacket
	);

	SoC_addr_router_002 addr_router_002 (
		.sink_ready         (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                    //          .valid
		.src_data           (addr_router_002_src_data),                                                     //          .data
		.src_channel        (addr_router_002_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                               //          .endofpacket
	);

	SoC_addr_router_003 addr_router_003 (
		.sink_ready         (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                           //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                           //          .valid
		.src_data           (addr_router_003_src_data),                                                            //          .data
		.src_channel        (addr_router_003_src_channel),                                                         //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                      //          .endofpacket
	);

	SoC_id_router id_router (
		.sink_ready         (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                               //       src.ready
		.src_valid          (id_router_src_valid),                                                               //          .valid
		.src_data           (id_router_src_data),                                                                //          .data
		.src_channel        (id_router_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                          //          .endofpacket
	);

	SoC_id_router id_router_001 (
		.sink_ready         (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ins_mem0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                //       src.ready
		.src_valid          (id_router_001_src_valid),                                                //          .valid
		.src_data           (id_router_001_src_data),                                                 //          .data
		.src_channel        (id_router_001_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                           //          .endofpacket
	);

	SoC_id_router id_router_002 (
		.sink_ready         (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_mem0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                 //       src.ready
		.src_valid          (id_router_002_src_valid),                                                 //          .valid
		.src_data           (id_router_002_src_data),                                                  //          .data
		.src_channel        (id_router_002_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                            //          .endofpacket
	);

	SoC_id_router id_router_003 (
		.sink_ready         (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                              //       src.ready
		.src_valid          (id_router_003_src_valid),                                              //          .valid
		.src_data           (id_router_003_src_data),                                               //          .data
		.src_channel        (id_router_003_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router id_router_004 (
		.sink_ready         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                  //       src.ready
		.src_valid          (id_router_004_src_valid),                                                  //          .valid
		.src_data           (id_router_004_src_data),                                                   //          .data
		.src_channel        (id_router_004_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_005 id_router_005 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                  //          .valid
		.src_data           (id_router_005_src_data),                                                                   //          .data
		.src_channel        (id_router_005_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_005 id_router_006 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                               //       src.ready
		.src_valid          (id_router_006_src_valid),                                               //          .valid
		.src_data           (id_router_006_src_data),                                                //          .data
		.src_channel        (id_router_006_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_007 id_router_007 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                        //       src.ready
		.src_valid          (id_router_007_src_valid),                                                        //          .valid
		.src_data           (id_router_007_src_data),                                                         //          .data
		.src_channel        (id_router_007_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                   //          .endofpacket
	);

	SoC_id_router_008 id_router_008 (
		.sink_ready         (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                           //       src.ready
		.src_valid          (id_router_008_src_valid),                                                           //          .valid
		.src_data           (id_router_008_src_data),                                                            //          .data
		.src_channel        (id_router_008_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                      //          .endofpacket
	);

	SoC_id_router_008 id_router_009 (
		.sink_ready         (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ins_mem1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                //       src.ready
		.src_valid          (id_router_009_src_valid),                                                //          .valid
		.src_data           (id_router_009_src_data),                                                 //          .data
		.src_channel        (id_router_009_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                           //          .endofpacket
	);

	SoC_id_router_010 id_router_010 (
		.sink_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_010_src_valid),                                                                  //          .valid
		.src_data           (id_router_010_src_data),                                                                   //          .data
		.src_channel        (id_router_010_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_010 id_router_011 (
		.sink_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                               //       src.ready
		.src_valid          (id_router_011_src_valid),                                               //          .valid
		.src_data           (id_router_011_src_data),                                                //          .data
		.src_channel        (id_router_011_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_008 id_router_012 (
		.sink_ready         (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                               //       src.ready
		.src_valid          (id_router_012_src_valid),                                               //          .valid
		.src_data           (id_router_012_src_data),                                                //          .data
		.src_channel        (id_router_012_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_008 id_router_013 (
		.sink_ready         (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_mem1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                 //       src.ready
		.src_valid          (id_router_013_src_valid),                                                 //          .valid
		.src_data           (id_router_013_src_data),                                                  //          .data
		.src_channel        (id_router_013_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                            //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (14),
		.VALID_WIDTH               (14),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),              //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),              //          .valid
		.cmd_sink_data          (addr_router_src_data),               //          .data
		.cmd_sink_channel       (addr_router_src_channel),            //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),             //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),             //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),           //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),              //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),     //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),       //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (14),
		.VALID_WIDTH               (14),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_003_src_data),           //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_003_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_003_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_003_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_003_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_003_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (cpu0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (cpu1_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (cpu1_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu0_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	SoC_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                            //        clk.clk
		.reset              (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),            //           .channel
		.sink_data          (limiter_cmd_src_data),               //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),    //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),          //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),          //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),           //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),        //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket)     //           .endofpacket
	);

	SoC_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //      src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //      src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_002_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_002_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_002_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_002_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_002_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_002_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_002_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_002_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_002_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_002_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_002_src5_endofpacket),   //          .endofpacket
		.src6_ready         (cmd_xbar_demux_002_src6_ready),         //      src6.ready
		.src6_valid         (cmd_xbar_demux_002_src6_valid),         //          .valid
		.src6_data          (cmd_xbar_demux_002_src6_data),          //          .data
		.src6_channel       (cmd_xbar_demux_002_src6_channel),       //          .channel
		.src6_startofpacket (cmd_xbar_demux_002_src6_startofpacket), //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_002_src6_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_003_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_003_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_003_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_003_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_003_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_003_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_003_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_003_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_003_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_003_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_003_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_003_src3_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_007 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src7_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_008 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src1_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_009 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src2_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_012 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_012_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_012_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_012_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_012_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_012_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_012_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src5_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src5_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src5_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src5_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src5_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src5_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src2_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_013 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_013_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_013_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_013_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_013_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_013_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_013_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src6_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src6_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src6_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src6_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src6_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src6_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_005 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_005 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_005 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_005 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_012_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_012_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_013_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_013_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_007_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_008_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_009_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_010_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_011_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_012_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_013_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_003 rsp_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_008_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_009_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_012_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_012_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_013_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_013_src1_endofpacket)    //          .endofpacket
	);

	SoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (cpu0_d_irq_irq)                      //    sender.irq
	);

	SoC_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (cpu1_d_irq_irq)                      //    sender.irq
	);

endmodule
