// SoC.v

// Generated using ACDS version 12.1 177 at 2022.02.25.14:55:15

`timescale 1 ps / 1 ps
module SoC (
		output wire [7:0]  led_out_external_connection_export, // led_out_external_connection.export
		output wire        pll_c2_clk,                         //                      pll_c2.clk
		output wire [12:0] sdram_control_wire_addr,            //          sdram_control_wire.addr
		output wire [1:0]  sdram_control_wire_ba,              //                            .ba
		output wire        sdram_control_wire_cas_n,           //                            .cas_n
		output wire        sdram_control_wire_cke,             //                            .cke
		output wire        sdram_control_wire_cs_n,            //                            .cs_n
		inout  wire [31:0] sdram_control_wire_dq,              //                            .dq
		output wire [3:0]  sdram_control_wire_dqm,             //                            .dqm
		output wire        sdram_control_wire_ras_n,           //                            .ras_n
		output wire        sdram_control_wire_we_n,            //                            .we_n
		input  wire        reset_reset_n,                      //                       reset.reset_n
		input  wire        clk_clk                             //                         clk.clk
	);

	wire          pll_c0_clk;                                                                                         // PLL:c0 -> [CRC_Custom_Instruction_0:clk, addr_router:clk, addr_router_001:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cpu:clk, cpu_data_master_translator:clk, cpu_data_master_translator_avalon_universal_master_0_agent:clk, cpu_instruction_master_translator:clk, cpu_instruction_master_translator_avalon_universal_master_0_agent:clk, cpu_jtag_debug_module_translator:clk, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, crosser:in_clk, crosser_001:out_clk, id_router:clk, id_router_001:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, led_out:clk, led_out_s1_translator:clk, led_out_s1_translator_avalon_universal_slave_0_agent:clk, led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, mm_clock_crossing_bridge_0:s0_clk, mm_clock_crossing_bridge_0_s0_translator:clk, mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:clk, mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller_001:clk, sdram_control:clk, sdram_control_s1_translator:clk, sdram_control_s1_translator_avalon_universal_slave_0_agent:clk, sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire          pll_c1_clk;                                                                                         // PLL:c1 -> [addr_router_002:clk, cmd_xbar_demux_002:clk, high_freq_timer:clk, high_freq_timer_s1_translator:clk, high_freq_timer_s1_translator_avalon_universal_slave_0_agent:clk, high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, limiter_001:clk, mm_clock_crossing_bridge_0:m0_clk, mm_clock_crossing_bridge_0_m0_translator:clk, mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_mux_002:clk, rst_controller_002:clk, sysid:clock, sysid_control_slave_translator:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer:clk, timer_s1_translator:clk, timer_s1_translator_avalon_universal_slave_0_agent:clk, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire   [31:0] cpu_custom_instruction_master_result;                                                               // cpu_custom_instruction_master_translator:ci_slave_result -> cpu:E_ci_combo_result
	wire    [4:0] cpu_custom_instruction_master_b;                                                                    // cpu:E_ci_combo_b -> cpu_custom_instruction_master_translator:ci_slave_b
	wire    [4:0] cpu_custom_instruction_master_c;                                                                    // cpu:E_ci_combo_c -> cpu_custom_instruction_master_translator:ci_slave_c
	wire   [31:0] cpu_custom_instruction_master_dataa;                                                                // cpu:E_ci_combo_dataa -> cpu_custom_instruction_master_translator:ci_slave_dataa
	wire    [4:0] cpu_custom_instruction_master_a;                                                                    // cpu:E_ci_combo_a -> cpu_custom_instruction_master_translator:ci_slave_a
	wire          cpu_custom_instruction_master_readra;                                                               // cpu:E_ci_combo_readra -> cpu_custom_instruction_master_translator:ci_slave_readra
	wire    [7:0] cpu_custom_instruction_master_n;                                                                    // cpu:E_ci_combo_n -> cpu_custom_instruction_master_translator:ci_slave_n
	wire          cpu_custom_instruction_master_writerc;                                                              // cpu:E_ci_combo_writerc -> cpu_custom_instruction_master_translator:ci_slave_writerc
	wire   [31:0] cpu_custom_instruction_master_datab;                                                                // cpu:E_ci_combo_datab -> cpu_custom_instruction_master_translator:ci_slave_datab
	wire          cpu_custom_instruction_master_readrb;                                                               // cpu:E_ci_combo_readrb -> cpu_custom_instruction_master_translator:ci_slave_readrb
	wire   [31:0] cpu_custom_instruction_master_ipending;                                                             // cpu:E_ci_combo_ipending -> cpu_custom_instruction_master_translator:ci_slave_ipending
	wire          cpu_custom_instruction_master_estatus;                                                              // cpu:E_ci_combo_estatus -> cpu_custom_instruction_master_translator:ci_slave_estatus
	wire   [31:0] cpu_custom_instruction_master_translator_comb_ci_master_result;                                     // cpu_custom_instruction_master_comb_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:comb_ci_master_result
	wire    [4:0] cpu_custom_instruction_master_translator_comb_ci_master_b;                                          // cpu_custom_instruction_master_translator:comb_ci_master_b -> cpu_custom_instruction_master_comb_xconnect:ci_slave_b
	wire    [4:0] cpu_custom_instruction_master_translator_comb_ci_master_c;                                          // cpu_custom_instruction_master_translator:comb_ci_master_c -> cpu_custom_instruction_master_comb_xconnect:ci_slave_c
	wire   [31:0] cpu_custom_instruction_master_translator_comb_ci_master_dataa;                                      // cpu_custom_instruction_master_translator:comb_ci_master_dataa -> cpu_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire    [4:0] cpu_custom_instruction_master_translator_comb_ci_master_a;                                          // cpu_custom_instruction_master_translator:comb_ci_master_a -> cpu_custom_instruction_master_comb_xconnect:ci_slave_a
	wire          cpu_custom_instruction_master_translator_comb_ci_master_readra;                                     // cpu_custom_instruction_master_translator:comb_ci_master_readra -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire    [7:0] cpu_custom_instruction_master_translator_comb_ci_master_n;                                          // cpu_custom_instruction_master_translator:comb_ci_master_n -> cpu_custom_instruction_master_comb_xconnect:ci_slave_n
	wire          cpu_custom_instruction_master_translator_comb_ci_master_writerc;                                    // cpu_custom_instruction_master_translator:comb_ci_master_writerc -> cpu_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [31:0] cpu_custom_instruction_master_translator_comb_ci_master_datab;                                      // cpu_custom_instruction_master_translator:comb_ci_master_datab -> cpu_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire   [31:0] cpu_custom_instruction_master_translator_comb_ci_master_ipending;                                   // cpu_custom_instruction_master_translator:comb_ci_master_ipending -> cpu_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire          cpu_custom_instruction_master_translator_comb_ci_master_readrb;                                     // cpu_custom_instruction_master_translator:comb_ci_master_readrb -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire          cpu_custom_instruction_master_translator_comb_ci_master_estatus;                                    // cpu_custom_instruction_master_translator:comb_ci_master_estatus -> cpu_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire   [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_result;                                      // cpu_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_comb_xconnect:ci_master0_result
	wire    [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_b;                                           // cpu_custom_instruction_master_comb_xconnect:ci_master0_b -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire    [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_c;                                           // cpu_custom_instruction_master_comb_xconnect:ci_master0_c -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire   [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa;                                       // cpu_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire    [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_a;                                           // cpu_custom_instruction_master_comb_xconnect:ci_master0_a -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire          cpu_custom_instruction_master_comb_xconnect_ci_master0_readra;                                      // cpu_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire    [7:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_n;                                           // cpu_custom_instruction_master_comb_xconnect:ci_master0_n -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire          cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc;                                     // cpu_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_datab;                                       // cpu_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire   [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending;                                    // cpu_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire          cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb;                                      // cpu_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire          cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus;                                     // cpu_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire   [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_result;                              // CRC_Custom_Instruction_0:result -> cpu_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire   [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa;                               // cpu_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> CRC_Custom_Instruction_0:dataa
	wire    [2:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_n;                                   // cpu_custom_instruction_master_comb_slave_translator0:ci_master_n -> CRC_Custom_Instruction_0:n
	wire          cpu_instruction_master_waitrequest;                                                                 // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [27:0] cpu_instruction_master_address;                                                                     // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                        // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                    // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                                                               // cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	wire          cpu_data_master_waitrequest;                                                                        // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                          // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [27:0] cpu_data_master_address;                                                                            // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                              // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                               // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                           // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                        // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire    [3:0] cpu_data_master_byteenable;                                                                         // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                     // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                       // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                    // cpu_jtag_debug_module_translator:av_chipselect -> cpu:jtag_debug_module_select
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                         // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                      // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                 // cpu_jtag_debug_module_translator:av_begintransfer -> cpu:jtag_debug_module_begintransfer
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                   // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                    // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire          sdram_control_s1_translator_avalon_anti_slave_0_waitrequest;                                        // sdram_control:za_waitrequest -> sdram_control_s1_translator:av_waitrequest
	wire   [31:0] sdram_control_s1_translator_avalon_anti_slave_0_writedata;                                          // sdram_control_s1_translator:av_writedata -> sdram_control:az_data
	wire   [24:0] sdram_control_s1_translator_avalon_anti_slave_0_address;                                            // sdram_control_s1_translator:av_address -> sdram_control:az_addr
	wire          sdram_control_s1_translator_avalon_anti_slave_0_chipselect;                                         // sdram_control_s1_translator:av_chipselect -> sdram_control:az_cs
	wire          sdram_control_s1_translator_avalon_anti_slave_0_write;                                              // sdram_control_s1_translator:av_write -> sdram_control:az_wr_n
	wire          sdram_control_s1_translator_avalon_anti_slave_0_read;                                               // sdram_control_s1_translator:av_read -> sdram_control:az_rd_n
	wire   [31:0] sdram_control_s1_translator_avalon_anti_slave_0_readdata;                                           // sdram_control:za_data -> sdram_control_s1_translator:av_readdata
	wire          sdram_control_s1_translator_avalon_anti_slave_0_readdatavalid;                                      // sdram_control:za_valid -> sdram_control_s1_translator:av_readdatavalid
	wire    [3:0] sdram_control_s1_translator_avalon_anti_slave_0_byteenable;                                         // sdram_control_s1_translator:av_byteenable -> sdram_control:az_be_n
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_writedata;                                             // PLL_pll_slave_translator:av_writedata -> PLL:writedata
	wire    [1:0] pll_pll_slave_translator_avalon_anti_slave_0_address;                                               // PLL_pll_slave_translator:av_address -> PLL:address
	wire          pll_pll_slave_translator_avalon_anti_slave_0_write;                                                 // PLL_pll_slave_translator:av_write -> PLL:write
	wire          pll_pll_slave_translator_avalon_anti_slave_0_read;                                                  // PLL_pll_slave_translator:av_read -> PLL:read
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_readdata;                                              // PLL:readdata -> PLL_pll_slave_translator:av_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                             // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                               // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                 // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                              // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                   // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                    // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] led_out_s1_translator_avalon_anti_slave_0_writedata;                                                // led_out_s1_translator:av_writedata -> led_out:writedata
	wire    [1:0] led_out_s1_translator_avalon_anti_slave_0_address;                                                  // led_out_s1_translator:av_address -> led_out:address
	wire          led_out_s1_translator_avalon_anti_slave_0_chipselect;                                               // led_out_s1_translator:av_chipselect -> led_out:chipselect
	wire          led_out_s1_translator_avalon_anti_slave_0_write;                                                    // led_out_s1_translator:av_write -> led_out:write_n
	wire   [31:0] led_out_s1_translator_avalon_anti_slave_0_readdata;                                                 // led_out:readdata -> led_out_s1_translator:av_readdata
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_waitrequest;                           // mm_clock_crossing_bridge_0:s0_waitrequest -> mm_clock_crossing_bridge_0_s0_translator:av_waitrequest
	wire    [0:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_burstcount;                            // mm_clock_crossing_bridge_0_s0_translator:av_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_writedata;                             // mm_clock_crossing_bridge_0_s0_translator:av_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	wire    [9:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_address;                               // mm_clock_crossing_bridge_0_s0_translator:av_address -> mm_clock_crossing_bridge_0:s0_address
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_write;                                 // mm_clock_crossing_bridge_0_s0_translator:av_write -> mm_clock_crossing_bridge_0:s0_write
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_read;                                  // mm_clock_crossing_bridge_0_s0_translator:av_read -> mm_clock_crossing_bridge_0:s0_read
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdata;                              // mm_clock_crossing_bridge_0:s0_readdata -> mm_clock_crossing_bridge_0_s0_translator:av_readdata
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_debugaccess;                           // mm_clock_crossing_bridge_0_s0_translator:av_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdatavalid;                         // mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_clock_crossing_bridge_0_s0_translator:av_readdatavalid
	wire    [3:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_byteenable;                            // mm_clock_crossing_bridge_0_s0_translator:av_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	wire    [0:0] mm_clock_crossing_bridge_0_m0_burstcount;                                                           // mm_clock_crossing_bridge_0:m0_burstcount -> mm_clock_crossing_bridge_0_m0_translator:av_burstcount
	wire          mm_clock_crossing_bridge_0_m0_waitrequest;                                                          // mm_clock_crossing_bridge_0_m0_translator:av_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	wire    [9:0] mm_clock_crossing_bridge_0_m0_address;                                                              // mm_clock_crossing_bridge_0:m0_address -> mm_clock_crossing_bridge_0_m0_translator:av_address
	wire   [31:0] mm_clock_crossing_bridge_0_m0_writedata;                                                            // mm_clock_crossing_bridge_0:m0_writedata -> mm_clock_crossing_bridge_0_m0_translator:av_writedata
	wire          mm_clock_crossing_bridge_0_m0_write;                                                                // mm_clock_crossing_bridge_0:m0_write -> mm_clock_crossing_bridge_0_m0_translator:av_write
	wire          mm_clock_crossing_bridge_0_m0_read;                                                                 // mm_clock_crossing_bridge_0:m0_read -> mm_clock_crossing_bridge_0_m0_translator:av_read
	wire   [31:0] mm_clock_crossing_bridge_0_m0_readdata;                                                             // mm_clock_crossing_bridge_0_m0_translator:av_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	wire          mm_clock_crossing_bridge_0_m0_debugaccess;                                                          // mm_clock_crossing_bridge_0:m0_debugaccess -> mm_clock_crossing_bridge_0_m0_translator:av_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_0_m0_byteenable;                                                           // mm_clock_crossing_bridge_0:m0_byteenable -> mm_clock_crossing_bridge_0_m0_translator:av_byteenable
	wire          mm_clock_crossing_bridge_0_m0_readdatavalid;                                                        // mm_clock_crossing_bridge_0_m0_translator:av_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                  // timer_s1_translator:av_writedata -> timer:writedata
	wire    [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                    // timer_s1_translator:av_address -> timer:address
	wire          timer_s1_translator_avalon_anti_slave_0_chipselect;                                                 // timer_s1_translator:av_chipselect -> timer:chipselect
	wire          timer_s1_translator_avalon_anti_slave_0_write;                                                      // timer_s1_translator:av_write -> timer:write_n
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                   // timer:readdata -> timer_s1_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                         // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                        // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [15:0] high_freq_timer_s1_translator_avalon_anti_slave_0_writedata;                                        // high_freq_timer_s1_translator:av_writedata -> high_freq_timer:writedata
	wire    [2:0] high_freq_timer_s1_translator_avalon_anti_slave_0_address;                                          // high_freq_timer_s1_translator:av_address -> high_freq_timer:address
	wire          high_freq_timer_s1_translator_avalon_anti_slave_0_chipselect;                                       // high_freq_timer_s1_translator:av_chipselect -> high_freq_timer:chipselect
	wire          high_freq_timer_s1_translator_avalon_anti_slave_0_write;                                            // high_freq_timer_s1_translator:av_write -> high_freq_timer:write_n
	wire   [15:0] high_freq_timer_s1_translator_avalon_anti_slave_0_readdata;                                         // high_freq_timer:readdata -> high_freq_timer_s1_translator:av_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                            // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                             // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                              // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                   // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                  // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                   // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                               // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                            // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                             // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                          // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                   // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                    // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                     // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_data_master_translator_avalon_universal_master_0_address;                                       // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                          // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                         // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                          // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                      // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                   // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                    // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                 // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [27:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                        // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // sdram_control_s1_translator:uav_waitrequest -> sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_control_s1_translator:uav_burstcount
	wire   [31:0] sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_control_s1_translator:uav_writedata
	wire   [27:0] sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_control_s1_translator:uav_address
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_control_s1_translator:uav_write
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_control_s1_translator:uav_lock
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_control_s1_translator:uav_read
	wire   [31:0] sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // sdram_control_s1_translator:uav_readdata -> sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // sdram_control_s1_translator:uav_readdatavalid -> sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_control_s1_translator:uav_debugaccess
	wire    [3:0] sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // sdram_control_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_control_s1_translator:uav_byteenable
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // sdram_control_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // sdram_control_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_control_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sdram_control_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // sdram_control_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_control_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // sdram_control_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_control_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // PLL_pll_slave_translator:uav_waitrequest -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> PLL_pll_slave_translator:uav_burstcount
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                               // PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> PLL_pll_slave_translator:uav_writedata
	wire   [27:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                                 // PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> PLL_pll_slave_translator:uav_address
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                                   // PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> PLL_pll_slave_translator:uav_write
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                    // PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> PLL_pll_slave_translator:uav_lock
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                                    // PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> PLL_pll_slave_translator:uav_read
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                // PLL_pll_slave_translator:uav_readdata -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // PLL_pll_slave_translator:uav_readdatavalid -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PLL_pll_slave_translator:uav_debugaccess
	wire    [3:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // PLL_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> PLL_pll_slave_translator:uav_byteenable
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                             // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PLL_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PLL_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // PLL_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                       // PLL_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                        // PLL_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                       // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PLL_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [27:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                  // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // led_out_s1_translator:uav_waitrequest -> led_out_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // led_out_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_out_s1_translator:uav_burstcount
	wire   [31:0] led_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // led_out_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_out_s1_translator:uav_writedata
	wire   [27:0] led_out_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // led_out_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_out_s1_translator:uav_address
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // led_out_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_out_s1_translator:uav_write
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // led_out_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_out_s1_translator:uav_lock
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // led_out_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_out_s1_translator:uav_read
	wire   [31:0] led_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // led_out_s1_translator:uav_readdata -> led_out_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // led_out_s1_translator:uav_readdatavalid -> led_out_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // led_out_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_out_s1_translator:uav_debugaccess
	wire    [3:0] led_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // led_out_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_out_s1_translator:uav_byteenable
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // led_out_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // led_out_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // led_out_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // led_out_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_out_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // led_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // led_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] led_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // led_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // led_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // mm_clock_crossing_bridge_0_s0_translator:uav_waitrequest -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> mm_clock_crossing_bridge_0_s0_translator:uav_burstcount
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata;               // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> mm_clock_crossing_bridge_0_s0_translator:uav_writedata
	wire   [27:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_address;                 // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> mm_clock_crossing_bridge_0_s0_translator:uav_address
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_write;                   // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> mm_clock_crossing_bridge_0_s0_translator:uav_write
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_lock;                    // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> mm_clock_crossing_bridge_0_s0_translator:uav_lock
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_read;                    // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> mm_clock_crossing_bridge_0_s0_translator:uav_read
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                // mm_clock_crossing_bridge_0_s0_translator:uav_readdata -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // mm_clock_crossing_bridge_0_s0_translator:uav_readdatavalid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mm_clock_crossing_bridge_0_s0_translator:uav_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> mm_clock_crossing_bridge_0_s0_translator:uav_byteenable
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data;             // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_waitrequest;                     // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> mm_clock_crossing_bridge_0_m0_translator:uav_waitrequest
	wire    [2:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_burstcount;                      // mm_clock_crossing_bridge_0_m0_translator:uav_burstcount -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_writedata;                       // mm_clock_crossing_bridge_0_m0_translator:uav_writedata -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire    [9:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_address;                         // mm_clock_crossing_bridge_0_m0_translator:uav_address -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_address
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_lock;                            // mm_clock_crossing_bridge_0_m0_translator:uav_lock -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_write;                           // mm_clock_crossing_bridge_0_m0_translator:uav_write -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_write
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_read;                            // mm_clock_crossing_bridge_0_m0_translator:uav_read -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdata;                        // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_readdata -> mm_clock_crossing_bridge_0_m0_translator:uav_readdata
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_debugaccess;                     // mm_clock_crossing_bridge_0_m0_translator:uav_debugaccess -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_byteenable;                      // mm_clock_crossing_bridge_0_m0_translator:uav_byteenable -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdatavalid;                   // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> mm_clock_crossing_bridge_0_m0_translator:uav_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire    [9:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire    [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire    [9:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // high_freq_timer_s1_translator:uav_waitrequest -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_freq_timer_s1_translator:uav_burstcount
	wire   [31:0] high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_freq_timer_s1_translator:uav_writedata
	wire    [9:0] high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_freq_timer_s1_translator:uav_address
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_freq_timer_s1_translator:uav_write
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_freq_timer_s1_translator:uav_lock
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_freq_timer_s1_translator:uav_read
	wire   [31:0] high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // high_freq_timer_s1_translator:uav_readdata -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // high_freq_timer_s1_translator:uav_readdatavalid -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_freq_timer_s1_translator:uav_debugaccess
	wire    [3:0] high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_freq_timer_s1_translator:uav_byteenable
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                         // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [100:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                          // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                          // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                        // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [100:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                 // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                // addr_router_001:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [100:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // sdram_control_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // sdram_control_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // sdram_control_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [100:0] sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // sdram_control_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_001:sink_ready -> sdram_control_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                   // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [100:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                                    // PLL_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_002:sink_ready -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [100:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_003:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // led_out_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // led_out_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // led_out_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [100:0] led_out_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // led_out_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          led_out_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_004:sink_ready -> led_out_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_valid;                   // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [100:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_data;                    // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;            // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_valid;                  // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;          // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [80:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_data;                   // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_ready;                  // addr_router_002:sink_ready -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [80:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_006:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [80:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_007:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [80:0] high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_008:sink_ready -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                        // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                              // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                      // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [100:0] addr_router_src_data;                                                                               // addr_router:src_data -> limiter:cmd_sink_data
	wire    [5:0] addr_router_src_channel;                                                                            // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                              // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                        // limiter:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                              // limiter:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                      // limiter:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [100:0] limiter_rsp_src_data;                                                                               // limiter:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_rsp_src_channel;                                                                            // limiter:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_002_src_endofpacket;                                                                    // addr_router_002:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_002_src_valid;                                                                          // addr_router_002:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_002_src_startofpacket;                                                                  // addr_router_002:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire   [80:0] addr_router_002_src_data;                                                                           // addr_router_002:src_data -> limiter_001:cmd_sink_data
	wire    [2:0] addr_router_002_src_channel;                                                                        // addr_router_002:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_002_src_ready;                                                                          // limiter_001:cmd_sink_ready -> addr_router_002:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                    // limiter_001:rsp_src_endofpacket -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                          // limiter_001:rsp_src_valid -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                  // limiter_001:rsp_src_startofpacket -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [80:0] limiter_001_rsp_src_data;                                                                           // limiter_001:rsp_src_data -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [2:0] limiter_001_rsp_src_channel;                                                                        // limiter_001:rsp_src_channel -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                          // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          rst_controller_reset_out_reset;                                                                     // rst_controller:reset_out -> [PLL:reset, PLL_pll_slave_translator:reset, PLL_pll_slave_translator_avalon_universal_slave_0_agent:reset, PLL_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, PLL_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_001:in_reset, id_router_002:reset, rsp_xbar_demux_002:reset]
	wire          cpu_jtag_debug_module_reset_reset;                                                                  // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire          rst_controller_001_reset_out_reset;                                                                 // rst_controller_001:reset_out -> [CRC_Custom_Instruction_0:reset, addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:out_reset, id_router:reset, id_router_001:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_out:reset_n, led_out_s1_translator:reset, led_out_s1_translator_avalon_universal_slave_0_agent:reset, led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, mm_clock_crossing_bridge_0:s0_reset, mm_clock_crossing_bridge_0_s0_translator:reset, mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:reset, mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram_control:reset_n, sdram_control_s1_translator:reset, sdram_control_s1_translator_avalon_universal_slave_0_agent:reset, sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_002_reset_out_reset;                                                                 // rst_controller_002:reset_out -> [addr_router_002:reset, cmd_xbar_demux_002:reset, high_freq_timer:reset_n, high_freq_timer_s1_translator:reset, high_freq_timer_s1_translator_avalon_universal_slave_0_agent:reset, high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, limiter_001:reset, mm_clock_crossing_bridge_0:m0_reset, mm_clock_crossing_bridge_0_m0_translator:reset, mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_mux_002:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                    // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                          // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                  // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [100:0] cmd_xbar_demux_src0_data;                                                                           // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [5:0] cmd_xbar_demux_src0_channel;                                                                        // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                          // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                    // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                          // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                  // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [100:0] cmd_xbar_demux_src1_data;                                                                           // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [5:0] cmd_xbar_demux_src1_channel;                                                                        // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                          // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                      // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                              // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src0_data;                                                                       // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [5:0] cmd_xbar_demux_001_src0_channel;                                                                    // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                      // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                      // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                              // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src1_data;                                                                       // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire    [5:0] cmd_xbar_demux_001_src1_channel;                                                                    // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                      // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                // cmd_xbar_demux_001:src3_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                      // cmd_xbar_demux_001:src3_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                              // cmd_xbar_demux_001:src3_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src3_data;                                                                       // cmd_xbar_demux_001:src3_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_demux_001_src3_channel;                                                                    // cmd_xbar_demux_001:src3_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                // cmd_xbar_demux_001:src4_endofpacket -> led_out_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                      // cmd_xbar_demux_001:src4_valid -> led_out_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                              // cmd_xbar_demux_001:src4_startofpacket -> led_out_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src4_data;                                                                       // cmd_xbar_demux_001:src4_data -> led_out_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_demux_001_src4_channel;                                                                    // cmd_xbar_demux_001:src4_channel -> led_out_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                // cmd_xbar_demux_001:src5_endofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                      // cmd_xbar_demux_001:src5_valid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                              // cmd_xbar_demux_001:src5_startofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src5_data;                                                                       // cmd_xbar_demux_001:src5_data -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_demux_001_src5_channel;                                                                    // cmd_xbar_demux_001:src5_channel -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                    // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                          // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                  // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [100:0] rsp_xbar_demux_src0_data;                                                                           // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [5:0] rsp_xbar_demux_src0_channel;                                                                        // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                          // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                    // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                          // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                  // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [100:0] rsp_xbar_demux_src1_data;                                                                           // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [5:0] rsp_xbar_demux_src1_channel;                                                                        // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                          // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                      // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                              // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [100:0] rsp_xbar_demux_001_src0_data;                                                                       // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [5:0] rsp_xbar_demux_001_src0_channel;                                                                    // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                      // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                      // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                              // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [100:0] rsp_xbar_demux_001_src1_data;                                                                       // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire    [5:0] rsp_xbar_demux_001_src1_channel;                                                                    // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                      // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                      // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                              // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [100:0] rsp_xbar_demux_003_src0_data;                                                                       // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire    [5:0] rsp_xbar_demux_003_src0_channel;                                                                    // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                      // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                      // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                              // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [100:0] rsp_xbar_demux_004_src0_data;                                                                       // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire    [5:0] rsp_xbar_demux_004_src0_channel;                                                                    // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                      // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                      // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                              // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [100:0] rsp_xbar_demux_005_src0_data;                                                                       // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire    [5:0] rsp_xbar_demux_005_src0_channel;                                                                    // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                      // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                        // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                      // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [100:0] limiter_cmd_src_data;                                                                               // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [5:0] limiter_cmd_src_channel;                                                                            // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                              // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                       // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                             // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                     // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [100:0] rsp_xbar_mux_src_data;                                                                              // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [5:0] rsp_xbar_mux_src_channel;                                                                           // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                             // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                    // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                          // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                  // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [100:0] addr_router_001_src_data;                                                                           // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [5:0] addr_router_001_src_channel;                                                                        // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                          // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                   // rsp_xbar_mux_001:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                         // rsp_xbar_mux_001:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                 // rsp_xbar_mux_001:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [100:0] rsp_xbar_mux_001_src_data;                                                                          // rsp_xbar_mux_001:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] rsp_xbar_mux_001_src_channel;                                                                       // rsp_xbar_mux_001:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                         // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                       // cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                             // cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                     // cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_mux_src_data;                                                                              // cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_src_channel;                                                                           // cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                          // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                        // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [100:0] id_router_src_data;                                                                                 // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [5:0] id_router_src_channel;                                                                              // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                   // cmd_xbar_mux_001:src_endofpacket -> sdram_control_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                         // cmd_xbar_mux_001:src_valid -> sdram_control_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                 // cmd_xbar_mux_001:src_startofpacket -> sdram_control_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_mux_001_src_data;                                                                          // cmd_xbar_mux_001:src_data -> sdram_control_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_001_src_channel;                                                                       // cmd_xbar_mux_001:src_channel -> sdram_control_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                         // sdram_control_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                      // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                            // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                    // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [100:0] id_router_001_src_data;                                                                             // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [5:0] id_router_001_src_channel;                                                                          // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          crosser_out_ready;                                                                                  // PLL_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_002_src_endofpacket;                                                                      // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                            // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                    // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [100:0] id_router_002_src_data;                                                                             // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [5:0] id_router_002_src_channel;                                                                          // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_003_src_endofpacket;                                                                      // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                            // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                    // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [100:0] id_router_003_src_data;                                                                             // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [5:0] id_router_003_src_channel;                                                                          // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                      // led_out_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                      // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                            // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                    // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [100:0] id_router_004_src_data;                                                                             // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [5:0] id_router_004_src_channel;                                                                          // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                      // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                      // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                            // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                    // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [100:0] id_router_005_src_data;                                                                             // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire    [5:0] id_router_005_src_channel;                                                                          // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                            // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                // cmd_xbar_demux_002:src0_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                      // cmd_xbar_demux_002:src0_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                              // cmd_xbar_demux_002:src0_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] cmd_xbar_demux_002_src0_data;                                                                       // cmd_xbar_demux_002:src0_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_002_src0_channel;                                                                    // cmd_xbar_demux_002:src0_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                                // cmd_xbar_demux_002:src1_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                      // cmd_xbar_demux_002:src1_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                              // cmd_xbar_demux_002:src1_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] cmd_xbar_demux_002_src1_data;                                                                       // cmd_xbar_demux_002:src1_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_002_src1_channel;                                                                    // cmd_xbar_demux_002:src1_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src2_endofpacket;                                                                // cmd_xbar_demux_002:src2_endofpacket -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src2_valid;                                                                      // cmd_xbar_demux_002:src2_valid -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src2_startofpacket;                                                              // cmd_xbar_demux_002:src2_startofpacket -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] cmd_xbar_demux_002_src2_data;                                                                       // cmd_xbar_demux_002:src2_data -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_002_src2_channel;                                                                    // cmd_xbar_demux_002:src2_channel -> high_freq_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                      // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                              // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire   [80:0] rsp_xbar_demux_006_src0_data;                                                                       // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_002:sink0_data
	wire    [2:0] rsp_xbar_demux_006_src0_channel;                                                                    // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                      // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                      // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_002:sink1_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                              // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire   [80:0] rsp_xbar_demux_007_src0_data;                                                                       // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_002:sink1_data
	wire    [2:0] rsp_xbar_demux_007_src0_channel;                                                                    // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_002:sink1_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                      // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                      // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_002:sink2_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                              // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire   [80:0] rsp_xbar_demux_008_src0_data;                                                                       // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_002:sink2_data
	wire    [2:0] rsp_xbar_demux_008_src0_channel;                                                                    // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_002:sink2_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                      // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_008:src0_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                    // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                  // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [80:0] limiter_001_cmd_src_data;                                                                           // limiter_001:cmd_src_data -> cmd_xbar_demux_002:sink_data
	wire    [2:0] limiter_001_cmd_src_channel;                                                                        // limiter_001:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                          // cmd_xbar_demux_002:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                   // rsp_xbar_mux_002:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                         // rsp_xbar_mux_002:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                                 // rsp_xbar_mux_002:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire   [80:0] rsp_xbar_mux_002_src_data;                                                                          // rsp_xbar_mux_002:src_data -> limiter_001:rsp_sink_data
	wire    [2:0] rsp_xbar_mux_002_src_channel;                                                                       // rsp_xbar_mux_002:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                         // limiter_001:rsp_sink_ready -> rsp_xbar_mux_002:src_ready
	wire          cmd_xbar_demux_002_src0_ready;                                                                      // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src0_ready
	wire          id_router_006_src_endofpacket;                                                                      // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                            // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                    // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [80:0] id_router_006_src_data;                                                                             // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire    [2:0] id_router_006_src_channel;                                                                          // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                            // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_002_src1_ready;                                                                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src1_ready
	wire          id_router_007_src_endofpacket;                                                                      // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                            // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                    // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [80:0] id_router_007_src_data;                                                                             // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire    [2:0] id_router_007_src_channel;                                                                          // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                            // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_002_src2_ready;                                                                      // high_freq_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src2_ready
	wire          id_router_008_src_endofpacket;                                                                      // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                            // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                    // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [80:0] id_router_008_src_data;                                                                             // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire    [2:0] id_router_008_src_channel;                                                                          // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                            // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          crosser_out_endofpacket;                                                                            // crosser:out_endofpacket -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                  // crosser:out_valid -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                          // crosser:out_startofpacket -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] crosser_out_data;                                                                                   // crosser:out_data -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] crosser_out_channel;                                                                                // crosser:out_channel -> PLL_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                // cmd_xbar_demux_001:src2_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                      // cmd_xbar_demux_001:src2_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                              // cmd_xbar_demux_001:src2_startofpacket -> crosser:in_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src2_data;                                                                       // cmd_xbar_demux_001:src2_data -> crosser:in_data
	wire    [5:0] cmd_xbar_demux_001_src2_channel;                                                                    // cmd_xbar_demux_001:src2_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                      // crosser:in_ready -> cmd_xbar_demux_001:src2_ready
	wire          crosser_001_out_endofpacket;                                                                        // crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          crosser_001_out_valid;                                                                              // crosser_001:out_valid -> rsp_xbar_mux_001:sink2_valid
	wire          crosser_001_out_startofpacket;                                                                      // crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [100:0] crosser_001_out_data;                                                                               // crosser_001:out_data -> rsp_xbar_mux_001:sink2_data
	wire    [5:0] crosser_001_out_channel;                                                                            // crosser_001:out_channel -> rsp_xbar_mux_001:sink2_channel
	wire          crosser_001_out_ready;                                                                              // rsp_xbar_mux_001:sink2_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                // rsp_xbar_demux_002:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                      // rsp_xbar_demux_002:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                              // rsp_xbar_demux_002:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [100:0] rsp_xbar_demux_002_src0_data;                                                                       // rsp_xbar_demux_002:src0_data -> crosser_001:in_data
	wire    [5:0] rsp_xbar_demux_002_src0_channel;                                                                    // rsp_xbar_demux_002:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                      // crosser_001:in_ready -> rsp_xbar_demux_002:src0_ready
	wire    [5:0] limiter_cmd_valid_data;                                                                             // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire    [2:0] limiter_001_cmd_valid_data;                                                                         // limiter_001:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	wire          irq_mapper_receiver1_irq;                                                                           // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                      // irq_mapper:sender_irq -> cpu:d_irq
	wire          irq_mapper_receiver0_irq;                                                                           // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                      // timer:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver2_irq;                                                                           // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                  // high_freq_timer:irq -> irq_synchronizer_001:receiver_irq

	SoC_PLL pll (
		.clk       (clk_clk),                                                //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                         // inclk_interface_reset.reset
		.read      (pll_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (pll_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (pll_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (pll_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (pll_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                             //                    c0.clk
		.c1        (pll_c1_clk),                                             //                    c1.clk
		.c2        (pll_c2_clk),                                             //                    c2.clk
		.areset    (),                                                       //        areset_conduit.export
		.locked    (),                                                       //        locked_conduit.export
		.phasedone ()                                                        //     phasedone_conduit.export
	);

	SoC_cpu cpu (
		.clk                                   (pll_c0_clk),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.E_ci_combo_result                     (cpu_custom_instruction_master_result),                               // custom_instruction_master.result
		.E_ci_combo_a                          (cpu_custom_instruction_master_a),                                    //                          .a
		.E_ci_combo_b                          (cpu_custom_instruction_master_b),                                    //                          .b
		.E_ci_combo_c                          (cpu_custom_instruction_master_c),                                    //                          .c
		.E_ci_combo_dataa                      (cpu_custom_instruction_master_dataa),                                //                          .dataa
		.E_ci_combo_datab                      (cpu_custom_instruction_master_datab),                                //                          .datab
		.E_ci_combo_estatus                    (cpu_custom_instruction_master_estatus),                              //                          .estatus
		.E_ci_combo_ipending                   (cpu_custom_instruction_master_ipending),                             //                          .ipending
		.E_ci_combo_n                          (cpu_custom_instruction_master_n),                                    //                          .n
		.E_ci_combo_readra                     (cpu_custom_instruction_master_readra),                               //                          .readra
		.E_ci_combo_readrb                     (cpu_custom_instruction_master_readrb),                               //                          .readrb
		.E_ci_combo_writerc                    (cpu_custom_instruction_master_writerc)                               //                          .writerc
	);

	SoC_sdram_control sdram_control (
		.clk            (pll_c0_clk),                                                    //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                           // reset.reset_n
		.az_addr        (sdram_control_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_control_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_control_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_control_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_control_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_control_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_control_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_control_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_control_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_control_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_control_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_control_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_control_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_control_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_control_wire_dq),                                         //      .export
		.zs_dqm         (sdram_control_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_control_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_control_wire_we_n)                                        //      .export
	);

	SoC_jtag_uart jtag_uart (
		.clk            (pll_c0_clk),                                                             //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                //               irq.irq
	);

	SoC_timer timer (
		.clk        (pll_c1_clk),                                         //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)                       //   irq.irq
	);

	SoC_sysid sysid (
		.clock    (pll_c1_clk),                                                  //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	SoC_led_out led_out (
		.clk        (pll_c0_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (led_out_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_out_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_out_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_out_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_out_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_out_external_connection_export)                    // external_connection.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_0 (
		.m0_clk           (pll_c1_clk),                                                                 //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                                         // m0_reset.reset
		.s0_clk           (pll_c0_clk),                                                                 //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                                         // s0_reset.reset
		.s0_waitrequest   (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_0_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_0_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_0_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_0_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_0_m0_writedata),                                    //         .writedata
		.m0_address       (mm_clock_crossing_bridge_0_m0_address),                                      //         .address
		.m0_write         (mm_clock_crossing_bridge_0_m0_write),                                        //         .write
		.m0_read          (mm_clock_crossing_bridge_0_m0_read),                                         //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_0_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_0_m0_debugaccess)                                   //         .debugaccess
	);

	SoC_high_freq_timer high_freq_timer (
		.clk        (pll_c1_clk),                                                   //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                          // reset.reset_n
		.address    (high_freq_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_freq_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_freq_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_freq_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_freq_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)                             //   irq.irq
	);

	CRC_Custom_Instruction #(
		.crc_width         (32),
		.polynomial_inital (34'b0011111111111111111111111111111111),
		.polynomial        (34'b0000000100110000010001110110110111),
		.reflected_input   (1),
		.reflected_output  (1),
		.xor_output        (34'b0011111111111111111111111111111111)
	) crc_custom_instruction_0 (
		.clk    (pll_c0_clk),                                                            //                         clock.clk
		.reset  (rst_controller_001_reset_out_reset),                                    //                         reset.reset
		.dataa  (cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.n      (cpu_custom_instruction_master_comb_slave_translator0_ci_master_n),      //                              .n
		.clk_en (),                                                                      //                              .clk_en
		.start  (),                                                                      //                              .start
		.done   (),                                                                      //                              .done
		.result (cpu_custom_instruction_master_comb_slave_translator0_ci_master_result)  //                              .result
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpu_custom_instruction_master_translator (
		.ci_slave_dataa          (cpu_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab          (cpu_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result         (cpu_custom_instruction_master_result),                             //               .result
		.ci_slave_n              (cpu_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra         (cpu_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb         (cpu_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc        (cpu_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a              (cpu_custom_instruction_master_a),                                  //               .a
		.ci_slave_b              (cpu_custom_instruction_master_b),                                  //               .b
		.ci_slave_c              (cpu_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending       (cpu_custom_instruction_master_ipending),                           //               .ipending
		.ci_slave_estatus        (cpu_custom_instruction_master_estatus),                            //               .estatus
		.comb_ci_master_dataa    (cpu_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab    (cpu_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result   (cpu_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n        (cpu_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra   (cpu_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb   (cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc  (cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a        (cpu_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b        (cpu_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c        (cpu_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending (cpu_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus  (cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk      (1'b0),                                                             //    (terminated)
		.ci_slave_multi_reset    (1'b0),                                                             //    (terminated)
		.ci_slave_multi_clken    (1'b0),                                                             //    (terminated)
		.ci_slave_multi_start    (1'b0),                                                             //    (terminated)
		.ci_slave_multi_done     (),                                                                 //    (terminated)
		.ci_slave_multi_dataa    (32'b00000000000000000000000000000000),                             //    (terminated)
		.ci_slave_multi_datab    (32'b00000000000000000000000000000000),                             //    (terminated)
		.ci_slave_multi_result   (),                                                                 //    (terminated)
		.ci_slave_multi_n        (8'b00000000),                                                      //    (terminated)
		.ci_slave_multi_readra   (1'b0),                                                             //    (terminated)
		.ci_slave_multi_readrb   (1'b0),                                                             //    (terminated)
		.ci_slave_multi_writerc  (1'b0),                                                             //    (terminated)
		.ci_slave_multi_a        (5'b00000),                                                         //    (terminated)
		.ci_slave_multi_b        (5'b00000),                                                         //    (terminated)
		.ci_slave_multi_c        (5'b00000),                                                         //    (terminated)
		.multi_ci_master_clk     (),                                                                 //    (terminated)
		.multi_ci_master_reset   (),                                                                 //    (terminated)
		.multi_ci_master_clken   (),                                                                 //    (terminated)
		.multi_ci_master_start   (),                                                                 //    (terminated)
		.multi_ci_master_done    (1'b0),                                                             //    (terminated)
		.multi_ci_master_dataa   (),                                                                 //    (terminated)
		.multi_ci_master_datab   (),                                                                 //    (terminated)
		.multi_ci_master_result  (32'b00000000000000000000000000000000),                             //    (terminated)
		.multi_ci_master_n       (),                                                                 //    (terminated)
		.multi_ci_master_readra  (),                                                                 //    (terminated)
		.multi_ci_master_readrb  (),                                                                 //    (terminated)
		.multi_ci_master_writerc (),                                                                 //    (terminated)
		.multi_ci_master_a       (),                                                                 //    (terminated)
		.multi_ci_master_b       (),                                                                 //    (terminated)
		.multi_ci_master_c       ()                                                                  //    (terminated)
	);

	SoC_cpu_custom_instruction_master_comb_xconnect cpu_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (cpu_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (cpu_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (cpu_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (cpu_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (cpu_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (cpu_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (cpu_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (cpu_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (cpu_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (cpu_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (cpu_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (cpu_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (cpu_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) cpu_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa     (cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab     (cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result    (cpu_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n         (cpu_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra    (cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb    (cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc   (cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a         (cpu_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b         (cpu_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c         (cpu_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending  (cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus   (cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa    (cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_result   (cpu_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n        (cpu_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_datab    (),                                                                      // (terminated)
		.ci_master_readra   (),                                                                      // (terminated)
		.ci_master_readrb   (),                                                                      // (terminated)
		.ci_master_writerc  (),                                                                      // (terminated)
		.ci_master_a        (),                                                                      // (terminated)
		.ci_master_b        (),                                                                      // (terminated)
		.ci_master_c        (),                                                                      // (terminated)
		.ci_master_ipending (),                                                                      // (terminated)
		.ci_master_estatus  (),                                                                      // (terminated)
		.ci_master_clk      (),                                                                      // (terminated)
		.ci_master_clken    (),                                                                      // (terminated)
		.ci_master_reset    (),                                                                      // (terminated)
		.ci_master_start    (),                                                                      // (terminated)
		.ci_master_done     (1'b0),                                                                  // (terminated)
		.ci_slave_clk       (1'b0),                                                                  // (terminated)
		.ci_slave_clken     (1'b0),                                                                  // (terminated)
		.ci_slave_reset     (1'b0),                                                                  // (terminated)
		.ci_slave_start     (1'b0),                                                                  // (terminated)
		.ci_slave_done      ()                                                                       // (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                   (pll_c0_clk),                                                                //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                        //                     reset.reset
		.uav_address           (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_write              (1'b0),                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                   (pll_c0_clk),                                                         //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_readdatavalid      (),                                                                   //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                   (pll_c0_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                               //                    reset.reset
		.uav_address           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_control_s1_translator (
		.clk                   (pll_c0_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address           (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_control_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_control_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_control_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_control_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_control_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_control_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_control_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_control_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_control_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pll_pll_slave_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pll_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pll_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pll_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pll_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pll_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (pll_c0_clk),                                                                             //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_out_s1_translator (
		.clk                   (pll_c0_clk),                                                            //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (led_out_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_out_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_out_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_out_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_out_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (led_out_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_out_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (led_out_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mm_clock_crossing_bridge_0_s0_translator (
		.clk                   (pll_c0_clk),                                                                               //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_chipselect         (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (10),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) mm_clock_crossing_bridge_0_m0_translator (
		.clk                   (pll_c1_clk),                                                                       //                       clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                               //                     reset.reset
		.uav_address           (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (mm_clock_crossing_bridge_0_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (mm_clock_crossing_bridge_0_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (mm_clock_crossing_bridge_0_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (mm_clock_crossing_bridge_0_m0_byteenable),                                         //                          .byteenable
		.av_read               (mm_clock_crossing_bridge_0_m0_read),                                               //                          .read
		.av_readdata           (mm_clock_crossing_bridge_0_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (mm_clock_crossing_bridge_0_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (mm_clock_crossing_bridge_0_m0_write),                                              //                          .write
		.av_writedata          (mm_clock_crossing_bridge_0_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (mm_clock_crossing_bridge_0_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                             //               (terminated)
		.av_begintransfer      (1'b0),                                                                             //               (terminated)
		.av_chipselect         (1'b0),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                             //               (terminated)
		.uav_clken             (),                                                                                 //               (terminated)
		.av_clken              (1'b1)                                                                              //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                   (pll_c1_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                  //                    reset.reset
		.uav_address           (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                   (pll_c1_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                             //                    reset.reset
		.uav_address           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_writedata          (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_freq_timer_s1_translator (
		.clk                   (pll_c1_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                            //                    reset.reset
		.uav_address           (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_freq_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_freq_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_freq_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_freq_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_freq_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (88),
		.PKT_THREAD_ID_H           (91),
		.PKT_THREAD_ID_L           (91),
		.PKT_CACHE_H               (98),
		.PKT_CACHE_L               (95),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_clk),                                                                         //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.av_address       (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                               //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (88),
		.PKT_THREAD_ID_H           (91),
		.PKT_THREAD_ID_L           (91),
		.PKT_CACHE_H               (98),
		.PKT_CACHE_L               (95),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_clk),                                                                  //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                  //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                   //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                          //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                            //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                   //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_control_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_control_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                          //                .channel
		.rf_sink_ready           (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_control_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_control_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_control_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_control_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_control_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_control_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_control_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_control_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                  //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                  //                .valid
		.cp_data                 (crosser_out_data),                                                                   //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                            //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                //                .channel
		.rf_sink_ready           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_out_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (led_out_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_out_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_out_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_out_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                 //                .channel
		.rf_sink_ready           (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                                    //                .channel
		.rf_sink_ready           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (9),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_BEGIN_BURST           (65),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.PKT_BURST_TYPE_H          (62),
		.PKT_BURST_TYPE_L          (61),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_TRANS_EXCLUSIVE       (51),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (69),
		.PKT_THREAD_ID_H           (71),
		.PKT_THREAD_ID_L           (71),
		.PKT_CACHE_H               (78),
		.PKT_CACHE_L               (75),
		.PKT_DATA_SIDEBAND_H       (64),
		.PKT_DATA_SIDEBAND_L       (64),
		.PKT_QOS_H                 (66),
		.PKT_QOS_L                 (66),
		.PKT_ADDR_SIDEBAND_H       (63),
		.PKT_ADDR_SIDEBAND_L       (63),
		.ST_DATA_W                 (81),
		.ST_CHANNEL_W              (3),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent (
		.clk              (pll_c1_clk),                                                                                //       clk.clk
		.reset            (rst_controller_002_reset_out_reset),                                                        // clk_reset.reset
		.av_address       (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                                 //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                                  //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                               //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                         //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                           //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                                  //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c1_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src0_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src0_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_002_src0_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src0_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src0_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src0_channel),                                               //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c1_clk),                                                                    //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c1_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src1_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src1_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_002_src1_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src1_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src1_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src1_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c1_clk),                                                                               //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_freq_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c1_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src2_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src2_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_002_src2_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src2_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src2_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src2_channel),                                                         //                .channel
		.rf_sink_ready           (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c1_clk),                                                                              //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	SoC_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_clk),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	SoC_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	SoC_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	SoC_id_router id_router_001 (
		.sink_ready         (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_control_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                     //       src.ready
		.src_valid          (id_router_001_src_valid),                                                     //          .valid
		.src_data           (id_router_001_src_data),                                                      //          .data
		.src_channel        (id_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                //          .endofpacket
	);

	SoC_id_router_002 id_router_002 (
		.sink_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                  //       src.ready
		.src_valid          (id_router_002_src_valid),                                                  //          .valid
		.src_data           (id_router_002_src_data),                                                   //          .data
		.src_channel        (id_router_002_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_002 id_router_003 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_clk),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                //          .valid
		.src_data           (id_router_003_src_data),                                                                 //          .data
		.src_channel        (id_router_003_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                           //          .endofpacket
	);

	SoC_id_router_002 id_router_004 (
		.sink_ready         (led_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_out_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                               //       src.ready
		.src_valid          (id_router_004_src_valid),                                               //          .valid
		.src_data           (id_router_004_src_data),                                                //          .data
		.src_channel        (id_router_004_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_002 id_router_005 (
		.sink_ready         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_clk),                                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                  //          .valid
		.src_data           (id_router_005_src_data),                                                                   //          .data
		.src_channel        (id_router_005_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_addr_router_002 addr_router_002 (
		.sink_ready         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c1_clk),                                                                                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                 //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                 //          .valid
		.src_data           (addr_router_002_src_data),                                                                  //          .data
		.src_channel        (addr_router_002_src_channel),                                                               //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                            //          .endofpacket
	);

	SoC_id_router_006 id_router_006 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c1_clk),                                                          //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                             //       src.ready
		.src_valid          (id_router_006_src_valid),                                             //          .valid
		.src_data           (id_router_006_src_data),                                              //          .data
		.src_channel        (id_router_006_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                        //          .endofpacket
	);

	SoC_id_router_006 id_router_007 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c1_clk),                                                                     //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                        //       src.ready
		.src_valid          (id_router_007_src_valid),                                                        //          .valid
		.src_data           (id_router_007_src_data),                                                         //          .data
		.src_channel        (id_router_007_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                   //          .endofpacket
	);

	SoC_id_router_006 id_router_008 (
		.sink_ready         (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_freq_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c1_clk),                                                                    //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                       //       src.ready
		.src_valid          (id_router_008_src_valid),                                                       //          .valid
		.src_data           (id_router_008_src_data),                                                        //          .data
		.src_channel        (id_router_008_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                  //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (88),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (pll_c0_clk),                         //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),              //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),              //          .valid
		.cmd_sink_data          (addr_router_src_data),               //          .data
		.cmd_sink_channel       (addr_router_src_channel),            //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),             //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),             //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),           //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),              //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),     //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),       //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (69),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (81),
		.ST_CHANNEL_W              (3),
		.VALID_WIDTH               (3),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (pll_c1_clk),                         //       clk.clk
		.reset                  (rst_controller_002_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_002_src_data),           //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_002_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_002_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_002_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_002_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_002_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                    // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                           //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_in2  (1'b0),                              // (terminated)
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (pll_c0_clk),                         //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (pll_c1_clk),                         //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	SoC_cmd_xbar_demux cmd_xbar_demux (
		.clk                (pll_c0_clk),                         //        clk.clk
		.reset              (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),            //           .channel
		.sink_data          (limiter_cmd_src_data),               //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)     //           .endofpacket
	);

	SoC_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (pll_c0_clk),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (pll_c0_clk),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (pll_c0_clk),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux (
		.clk                (pll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (pll_c0_clk),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (pll_c0_clk),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (pll_c0_clk),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (pll_c0_clk),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (pll_c0_clk),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (pll_c0_clk),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (crosser_001_out_ready),                 //     sink2.ready
		.sink2_valid         (crosser_001_out_valid),                 //          .valid
		.sink2_channel       (crosser_001_out_channel),               //          .channel
		.sink2_data          (crosser_001_out_data),                  //          .data
		.sink2_startofpacket (crosser_001_out_startofpacket),         //          .startofpacket
		.sink2_endofpacket   (crosser_001_out_endofpacket),           //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (pll_c1_clk),                            //        clk.clk
		.reset              (rst_controller_002_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_002_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_002_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_002_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_002_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket)    //           .endofpacket
	);

	SoC_rsp_xbar_demux_006 rsp_xbar_demux_006 (
		.clk                (pll_c1_clk),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_006 rsp_xbar_demux_007 (
		.clk                (pll_c1_clk),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_006 rsp_xbar_demux_008 (
		.clk                (pll_c1_clk),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (pll_c1_clk),                            //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_006_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_007_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_008_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (101),
		.BITS_PER_SYMBOL     (101),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (pll_c0_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src2_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src2_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src2_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src2_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src2_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (101),
		.BITS_PER_SYMBOL     (101),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (pll_c0_clk),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_002_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_002_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_002_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_002_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	SoC_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_c1_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_c1_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

endmodule
