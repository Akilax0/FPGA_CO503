// SoC.v

// Generated using ACDS version 12.1 177 at 2022.04.13.20:56:19

`timescale 1 ps / 1 ps
module SoC (
		input  wire  reset_reset_n, // reset.reset_n
		input  wire  clk_clk        //   clk.clk
	);

	wire         cpu_0_instruction_master_waitrequest;                                                               // cpu_0_instruction_master_translator:av_waitrequest -> cpu_0:i_waitrequest
	wire  [13:0] cpu_0_instruction_master_address;                                                                   // cpu_0:i_address -> cpu_0_instruction_master_translator:av_address
	wire         cpu_0_instruction_master_read;                                                                      // cpu_0:i_read -> cpu_0_instruction_master_translator:av_read
	wire  [31:0] cpu_0_instruction_master_readdata;                                                                  // cpu_0_instruction_master_translator:av_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_readdatavalid;                                                             // cpu_0_instruction_master_translator:av_readdatavalid -> cpu_0:i_readdatavalid
	wire         cpu_5_instruction_master_waitrequest;                                                               // cpu_5_instruction_master_translator:av_waitrequest -> cpu_5:i_waitrequest
	wire  [13:0] cpu_5_instruction_master_address;                                                                   // cpu_5:i_address -> cpu_5_instruction_master_translator:av_address
	wire         cpu_5_instruction_master_read;                                                                      // cpu_5:i_read -> cpu_5_instruction_master_translator:av_read
	wire  [31:0] cpu_5_instruction_master_readdata;                                                                  // cpu_5_instruction_master_translator:av_readdata -> cpu_5:i_readdata
	wire         cpu_5_instruction_master_readdatavalid;                                                             // cpu_5_instruction_master_translator:av_readdatavalid -> cpu_5:i_readdatavalid
	wire         cpu_5_data_master_waitrequest;                                                                      // cpu_5_data_master_translator:av_waitrequest -> cpu_5:d_waitrequest
	wire  [31:0] cpu_5_data_master_writedata;                                                                        // cpu_5:d_writedata -> cpu_5_data_master_translator:av_writedata
	wire  [13:0] cpu_5_data_master_address;                                                                          // cpu_5:d_address -> cpu_5_data_master_translator:av_address
	wire         cpu_5_data_master_write;                                                                            // cpu_5:d_write -> cpu_5_data_master_translator:av_write
	wire         cpu_5_data_master_read;                                                                             // cpu_5:d_read -> cpu_5_data_master_translator:av_read
	wire  [31:0] cpu_5_data_master_readdata;                                                                         // cpu_5_data_master_translator:av_readdata -> cpu_5:d_readdata
	wire         cpu_5_data_master_debugaccess;                                                                      // cpu_5:jtag_debug_module_debugaccess_to_roms -> cpu_5_data_master_translator:av_debugaccess
	wire   [3:0] cpu_5_data_master_byteenable;                                                                       // cpu_5:d_byteenable -> cpu_5_data_master_translator:av_byteenable
	wire         cpu_0_data_master_waitrequest;                                                                      // cpu_0_data_master_translator:av_waitrequest -> cpu_0:d_waitrequest
	wire  [31:0] cpu_0_data_master_writedata;                                                                        // cpu_0:d_writedata -> cpu_0_data_master_translator:av_writedata
	wire  [13:0] cpu_0_data_master_address;                                                                          // cpu_0:d_address -> cpu_0_data_master_translator:av_address
	wire         cpu_0_data_master_write;                                                                            // cpu_0:d_write -> cpu_0_data_master_translator:av_write
	wire         cpu_0_data_master_read;                                                                             // cpu_0:d_read -> cpu_0_data_master_translator:av_read
	wire  [31:0] cpu_0_data_master_readdata;                                                                         // cpu_0_data_master_translator:av_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_debugaccess;                                                                      // cpu_0:jtag_debug_module_debugaccess_to_roms -> cpu_0_data_master_translator:av_debugaccess
	wire   [3:0] cpu_0_data_master_byteenable;                                                                       // cpu_0:d_byteenable -> cpu_0_data_master_translator:av_byteenable
	wire         cpu_4_instruction_master_waitrequest;                                                               // cpu_4_instruction_master_translator:av_waitrequest -> cpu_4:i_waitrequest
	wire  [13:0] cpu_4_instruction_master_address;                                                                   // cpu_4:i_address -> cpu_4_instruction_master_translator:av_address
	wire         cpu_4_instruction_master_read;                                                                      // cpu_4:i_read -> cpu_4_instruction_master_translator:av_read
	wire  [31:0] cpu_4_instruction_master_readdata;                                                                  // cpu_4_instruction_master_translator:av_readdata -> cpu_4:i_readdata
	wire         cpu_4_instruction_master_readdatavalid;                                                             // cpu_4_instruction_master_translator:av_readdatavalid -> cpu_4:i_readdatavalid
	wire         cpu_4_data_master_waitrequest;                                                                      // cpu_4_data_master_translator:av_waitrequest -> cpu_4:d_waitrequest
	wire  [31:0] cpu_4_data_master_writedata;                                                                        // cpu_4:d_writedata -> cpu_4_data_master_translator:av_writedata
	wire  [13:0] cpu_4_data_master_address;                                                                          // cpu_4:d_address -> cpu_4_data_master_translator:av_address
	wire         cpu_4_data_master_write;                                                                            // cpu_4:d_write -> cpu_4_data_master_translator:av_write
	wire         cpu_4_data_master_read;                                                                             // cpu_4:d_read -> cpu_4_data_master_translator:av_read
	wire  [31:0] cpu_4_data_master_readdata;                                                                         // cpu_4_data_master_translator:av_readdata -> cpu_4:d_readdata
	wire         cpu_4_data_master_debugaccess;                                                                      // cpu_4:jtag_debug_module_debugaccess_to_roms -> cpu_4_data_master_translator:av_debugaccess
	wire   [3:0] cpu_4_data_master_byteenable;                                                                       // cpu_4:d_byteenable -> cpu_4_data_master_translator:av_byteenable
	wire         cpu_3_instruction_master_waitrequest;                                                               // cpu_3_instruction_master_translator:av_waitrequest -> cpu_3:i_waitrequest
	wire  [13:0] cpu_3_instruction_master_address;                                                                   // cpu_3:i_address -> cpu_3_instruction_master_translator:av_address
	wire         cpu_3_instruction_master_read;                                                                      // cpu_3:i_read -> cpu_3_instruction_master_translator:av_read
	wire  [31:0] cpu_3_instruction_master_readdata;                                                                  // cpu_3_instruction_master_translator:av_readdata -> cpu_3:i_readdata
	wire         cpu_3_instruction_master_readdatavalid;                                                             // cpu_3_instruction_master_translator:av_readdatavalid -> cpu_3:i_readdatavalid
	wire         cpu_3_data_master_waitrequest;                                                                      // cpu_3_data_master_translator:av_waitrequest -> cpu_3:d_waitrequest
	wire  [31:0] cpu_3_data_master_writedata;                                                                        // cpu_3:d_writedata -> cpu_3_data_master_translator:av_writedata
	wire  [13:0] cpu_3_data_master_address;                                                                          // cpu_3:d_address -> cpu_3_data_master_translator:av_address
	wire         cpu_3_data_master_write;                                                                            // cpu_3:d_write -> cpu_3_data_master_translator:av_write
	wire         cpu_3_data_master_read;                                                                             // cpu_3:d_read -> cpu_3_data_master_translator:av_read
	wire  [31:0] cpu_3_data_master_readdata;                                                                         // cpu_3_data_master_translator:av_readdata -> cpu_3:d_readdata
	wire         cpu_3_data_master_debugaccess;                                                                      // cpu_3:jtag_debug_module_debugaccess_to_roms -> cpu_3_data_master_translator:av_debugaccess
	wire   [3:0] cpu_3_data_master_byteenable;                                                                       // cpu_3:d_byteenable -> cpu_3_data_master_translator:av_byteenable
	wire         cpu_2_data_master_waitrequest;                                                                      // cpu_2_data_master_translator:av_waitrequest -> cpu_2:d_waitrequest
	wire  [31:0] cpu_2_data_master_writedata;                                                                        // cpu_2:d_writedata -> cpu_2_data_master_translator:av_writedata
	wire  [13:0] cpu_2_data_master_address;                                                                          // cpu_2:d_address -> cpu_2_data_master_translator:av_address
	wire         cpu_2_data_master_write;                                                                            // cpu_2:d_write -> cpu_2_data_master_translator:av_write
	wire         cpu_2_data_master_read;                                                                             // cpu_2:d_read -> cpu_2_data_master_translator:av_read
	wire  [31:0] cpu_2_data_master_readdata;                                                                         // cpu_2_data_master_translator:av_readdata -> cpu_2:d_readdata
	wire         cpu_2_data_master_debugaccess;                                                                      // cpu_2:jtag_debug_module_debugaccess_to_roms -> cpu_2_data_master_translator:av_debugaccess
	wire   [3:0] cpu_2_data_master_byteenable;                                                                       // cpu_2:d_byteenable -> cpu_2_data_master_translator:av_byteenable
	wire         cpu_2_instruction_master_waitrequest;                                                               // cpu_2_instruction_master_translator:av_waitrequest -> cpu_2:i_waitrequest
	wire  [13:0] cpu_2_instruction_master_address;                                                                   // cpu_2:i_address -> cpu_2_instruction_master_translator:av_address
	wire         cpu_2_instruction_master_read;                                                                      // cpu_2:i_read -> cpu_2_instruction_master_translator:av_read
	wire  [31:0] cpu_2_instruction_master_readdata;                                                                  // cpu_2_instruction_master_translator:av_readdata -> cpu_2:i_readdata
	wire         cpu_2_instruction_master_readdatavalid;                                                             // cpu_2_instruction_master_translator:av_readdatavalid -> cpu_2:i_readdatavalid
	wire         cpu_1_instruction_master_waitrequest;                                                               // cpu_1_instruction_master_translator:av_waitrequest -> cpu_1:i_waitrequest
	wire  [13:0] cpu_1_instruction_master_address;                                                                   // cpu_1:i_address -> cpu_1_instruction_master_translator:av_address
	wire         cpu_1_instruction_master_read;                                                                      // cpu_1:i_read -> cpu_1_instruction_master_translator:av_read
	wire  [31:0] cpu_1_instruction_master_readdata;                                                                  // cpu_1_instruction_master_translator:av_readdata -> cpu_1:i_readdata
	wire         cpu_1_instruction_master_readdatavalid;                                                             // cpu_1_instruction_master_translator:av_readdatavalid -> cpu_1:i_readdatavalid
	wire         cpu_1_data_master_waitrequest;                                                                      // cpu_1_data_master_translator:av_waitrequest -> cpu_1:d_waitrequest
	wire  [31:0] cpu_1_data_master_writedata;                                                                        // cpu_1:d_writedata -> cpu_1_data_master_translator:av_writedata
	wire  [13:0] cpu_1_data_master_address;                                                                          // cpu_1:d_address -> cpu_1_data_master_translator:av_address
	wire         cpu_1_data_master_write;                                                                            // cpu_1:d_write -> cpu_1_data_master_translator:av_write
	wire         cpu_1_data_master_read;                                                                             // cpu_1:d_read -> cpu_1_data_master_translator:av_read
	wire  [31:0] cpu_1_data_master_readdata;                                                                         // cpu_1_data_master_translator:av_readdata -> cpu_1:d_readdata
	wire         cpu_1_data_master_debugaccess;                                                                      // cpu_1:jtag_debug_module_debugaccess_to_roms -> cpu_1_data_master_translator:av_debugaccess
	wire   [3:0] cpu_1_data_master_byteenable;                                                                       // cpu_1:d_byteenable -> cpu_1_data_master_translator:av_byteenable
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_0_jtag_debug_module_translator:av_writedata -> cpu_0:jtag_debug_module_writedata
	wire   [8:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_0_jtag_debug_module_translator:av_address -> cpu_0:jtag_debug_module_address
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_0_jtag_debug_module_translator:av_chipselect -> cpu_0:jtag_debug_module_select
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_0_jtag_debug_module_translator:av_write -> cpu_0:jtag_debug_module_write
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_0:jtag_debug_module_readdata -> cpu_0_jtag_debug_module_translator:av_readdata
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_0_jtag_debug_module_translator:av_begintransfer -> cpu_0:jtag_debug_module_begintransfer
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_0_jtag_debug_module_translator:av_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire   [3:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_0_jtag_debug_module_translator:av_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire  [31:0] ins_mem_0_s1_translator_avalon_anti_slave_0_writedata;                                              // ins_mem_0_s1_translator:av_writedata -> ins_mem_0:writedata
	wire   [9:0] ins_mem_0_s1_translator_avalon_anti_slave_0_address;                                                // ins_mem_0_s1_translator:av_address -> ins_mem_0:address
	wire         ins_mem_0_s1_translator_avalon_anti_slave_0_chipselect;                                             // ins_mem_0_s1_translator:av_chipselect -> ins_mem_0:chipselect
	wire         ins_mem_0_s1_translator_avalon_anti_slave_0_clken;                                                  // ins_mem_0_s1_translator:av_clken -> ins_mem_0:clken
	wire         ins_mem_0_s1_translator_avalon_anti_slave_0_write;                                                  // ins_mem_0_s1_translator:av_write -> ins_mem_0:write
	wire  [31:0] ins_mem_0_s1_translator_avalon_anti_slave_0_readdata;                                               // ins_mem_0:readdata -> ins_mem_0_s1_translator:av_readdata
	wire   [3:0] ins_mem_0_s1_translator_avalon_anti_slave_0_byteenable;                                             // ins_mem_0_s1_translator:av_byteenable -> ins_mem_0:byteenable
	wire         atob_0_in_translator_avalon_anti_slave_0_waitrequest;                                               // atob_0:avalonmm_write_slave_waitrequest -> atob_0_in_translator:av_waitrequest
	wire  [31:0] atob_0_in_translator_avalon_anti_slave_0_writedata;                                                 // atob_0_in_translator:av_writedata -> atob_0:avalonmm_write_slave_writedata
	wire         atob_0_in_translator_avalon_anti_slave_0_write;                                                     // atob_0_in_translator:av_write -> atob_0:avalonmm_write_slave_write
	wire  [31:0] atob_0_in_csr_translator_avalon_anti_slave_0_writedata;                                             // atob_0_in_csr_translator:av_writedata -> atob_0:wrclk_control_slave_writedata
	wire   [2:0] atob_0_in_csr_translator_avalon_anti_slave_0_address;                                               // atob_0_in_csr_translator:av_address -> atob_0:wrclk_control_slave_address
	wire         atob_0_in_csr_translator_avalon_anti_slave_0_write;                                                 // atob_0_in_csr_translator:av_write -> atob_0:wrclk_control_slave_write
	wire         atob_0_in_csr_translator_avalon_anti_slave_0_read;                                                  // atob_0_in_csr_translator:av_read -> atob_0:wrclk_control_slave_read
	wire  [31:0] atob_0_in_csr_translator_avalon_anti_slave_0_readdata;                                              // atob_0:wrclk_control_slave_readdata -> atob_0_in_csr_translator:av_readdata
	wire         atob_0_out_translator_avalon_anti_slave_0_waitrequest;                                              // atob_0:avalonmm_read_slave_waitrequest -> atob_0_out_translator:av_waitrequest
	wire         atob_0_out_translator_avalon_anti_slave_0_read;                                                     // atob_0_out_translator:av_read -> atob_0:avalonmm_read_slave_read
	wire  [31:0] atob_0_out_translator_avalon_anti_slave_0_readdata;                                                 // atob_0:avalonmm_read_slave_readdata -> atob_0_out_translator:av_readdata
	wire         atob_1_in_translator_avalon_anti_slave_0_waitrequest;                                               // atob_1:avalonmm_write_slave_waitrequest -> atob_1_in_translator:av_waitrequest
	wire  [31:0] atob_1_in_translator_avalon_anti_slave_0_writedata;                                                 // atob_1_in_translator:av_writedata -> atob_1:avalonmm_write_slave_writedata
	wire         atob_1_in_translator_avalon_anti_slave_0_write;                                                     // atob_1_in_translator:av_write -> atob_1:avalonmm_write_slave_write
	wire  [31:0] atob_1_in_csr_translator_avalon_anti_slave_0_writedata;                                             // atob_1_in_csr_translator:av_writedata -> atob_1:wrclk_control_slave_writedata
	wire   [2:0] atob_1_in_csr_translator_avalon_anti_slave_0_address;                                               // atob_1_in_csr_translator:av_address -> atob_1:wrclk_control_slave_address
	wire         atob_1_in_csr_translator_avalon_anti_slave_0_write;                                                 // atob_1_in_csr_translator:av_write -> atob_1:wrclk_control_slave_write
	wire         atob_1_in_csr_translator_avalon_anti_slave_0_read;                                                  // atob_1_in_csr_translator:av_read -> atob_1:wrclk_control_slave_read
	wire  [31:0] atob_1_in_csr_translator_avalon_anti_slave_0_readdata;                                              // atob_1:wrclk_control_slave_readdata -> atob_1_in_csr_translator:av_readdata
	wire         atob_1_out_translator_avalon_anti_slave_0_waitrequest;                                              // atob_1:avalonmm_read_slave_waitrequest -> atob_1_out_translator:av_waitrequest
	wire         atob_1_out_translator_avalon_anti_slave_0_read;                                                     // atob_1_out_translator:av_read -> atob_1:avalonmm_read_slave_read
	wire  [31:0] atob_1_out_translator_avalon_anti_slave_0_readdata;                                                 // atob_1:avalonmm_read_slave_readdata -> atob_1_out_translator:av_readdata
	wire         atob_2_in_translator_avalon_anti_slave_0_waitrequest;                                               // atob_2:avalonmm_write_slave_waitrequest -> atob_2_in_translator:av_waitrequest
	wire  [31:0] atob_2_in_translator_avalon_anti_slave_0_writedata;                                                 // atob_2_in_translator:av_writedata -> atob_2:avalonmm_write_slave_writedata
	wire         atob_2_in_translator_avalon_anti_slave_0_write;                                                     // atob_2_in_translator:av_write -> atob_2:avalonmm_write_slave_write
	wire  [31:0] atob_2_in_csr_translator_avalon_anti_slave_0_writedata;                                             // atob_2_in_csr_translator:av_writedata -> atob_2:wrclk_control_slave_writedata
	wire   [2:0] atob_2_in_csr_translator_avalon_anti_slave_0_address;                                               // atob_2_in_csr_translator:av_address -> atob_2:wrclk_control_slave_address
	wire         atob_2_in_csr_translator_avalon_anti_slave_0_write;                                                 // atob_2_in_csr_translator:av_write -> atob_2:wrclk_control_slave_write
	wire         atob_2_in_csr_translator_avalon_anti_slave_0_read;                                                  // atob_2_in_csr_translator:av_read -> atob_2:wrclk_control_slave_read
	wire  [31:0] atob_2_in_csr_translator_avalon_anti_slave_0_readdata;                                              // atob_2:wrclk_control_slave_readdata -> atob_2_in_csr_translator:av_readdata
	wire         atob_2_out_translator_avalon_anti_slave_0_waitrequest;                                              // atob_2:avalonmm_read_slave_waitrequest -> atob_2_out_translator:av_waitrequest
	wire         atob_2_out_translator_avalon_anti_slave_0_read;                                                     // atob_2_out_translator:av_read -> atob_2:avalonmm_read_slave_read
	wire  [31:0] atob_2_out_translator_avalon_anti_slave_0_readdata;                                                 // atob_2:avalonmm_read_slave_readdata -> atob_2_out_translator:av_readdata
	wire         atod_0_in_translator_avalon_anti_slave_0_waitrequest;                                               // atod_0:avalonmm_write_slave_waitrequest -> atod_0_in_translator:av_waitrequest
	wire  [31:0] atod_0_in_translator_avalon_anti_slave_0_writedata;                                                 // atod_0_in_translator:av_writedata -> atod_0:avalonmm_write_slave_writedata
	wire         atod_0_in_translator_avalon_anti_slave_0_write;                                                     // atod_0_in_translator:av_write -> atod_0:avalonmm_write_slave_write
	wire         atod_0_out_translator_avalon_anti_slave_0_waitrequest;                                              // atod_0:avalonmm_read_slave_waitrequest -> atod_0_out_translator:av_waitrequest
	wire         atod_0_out_translator_avalon_anti_slave_0_read;                                                     // atod_0_out_translator:av_read -> atod_0:avalonmm_read_slave_read
	wire  [31:0] atod_0_out_translator_avalon_anti_slave_0_readdata;                                                 // atod_0:avalonmm_read_slave_readdata -> atod_0_out_translator:av_readdata
	wire  [31:0] atod_0_in_csr_translator_avalon_anti_slave_0_writedata;                                             // atod_0_in_csr_translator:av_writedata -> atod_0:wrclk_control_slave_writedata
	wire   [2:0] atod_0_in_csr_translator_avalon_anti_slave_0_address;                                               // atod_0_in_csr_translator:av_address -> atod_0:wrclk_control_slave_address
	wire         atod_0_in_csr_translator_avalon_anti_slave_0_write;                                                 // atod_0_in_csr_translator:av_write -> atod_0:wrclk_control_slave_write
	wire         atod_0_in_csr_translator_avalon_anti_slave_0_read;                                                  // atod_0_in_csr_translator:av_read -> atod_0:wrclk_control_slave_read
	wire  [31:0] atod_0_in_csr_translator_avalon_anti_slave_0_readdata;                                              // atod_0:wrclk_control_slave_readdata -> atod_0_in_csr_translator:av_readdata
	wire         atoe_0_in_translator_avalon_anti_slave_0_waitrequest;                                               // atoe_0:avalonmm_write_slave_waitrequest -> atoe_0_in_translator:av_waitrequest
	wire  [31:0] atoe_0_in_translator_avalon_anti_slave_0_writedata;                                                 // atoe_0_in_translator:av_writedata -> atoe_0:avalonmm_write_slave_writedata
	wire         atoe_0_in_translator_avalon_anti_slave_0_write;                                                     // atoe_0_in_translator:av_write -> atoe_0:avalonmm_write_slave_write
	wire         atoe_0_out_translator_avalon_anti_slave_0_waitrequest;                                              // atoe_0:avalonmm_read_slave_waitrequest -> atoe_0_out_translator:av_waitrequest
	wire         atoe_0_out_translator_avalon_anti_slave_0_read;                                                     // atoe_0_out_translator:av_read -> atoe_0:avalonmm_read_slave_read
	wire  [31:0] atoe_0_out_translator_avalon_anti_slave_0_readdata;                                                 // atoe_0:avalonmm_read_slave_readdata -> atoe_0_out_translator:av_readdata
	wire  [31:0] atoe_0_in_csr_translator_avalon_anti_slave_0_writedata;                                             // atoe_0_in_csr_translator:av_writedata -> atoe_0:wrclk_control_slave_writedata
	wire   [2:0] atoe_0_in_csr_translator_avalon_anti_slave_0_address;                                               // atoe_0_in_csr_translator:av_address -> atoe_0:wrclk_control_slave_address
	wire         atoe_0_in_csr_translator_avalon_anti_slave_0_write;                                                 // atoe_0_in_csr_translator:av_write -> atoe_0:wrclk_control_slave_write
	wire         atoe_0_in_csr_translator_avalon_anti_slave_0_read;                                                  // atoe_0_in_csr_translator:av_read -> atoe_0:wrclk_control_slave_read
	wire  [31:0] atoe_0_in_csr_translator_avalon_anti_slave_0_readdata;                                              // atoe_0:wrclk_control_slave_readdata -> atoe_0_in_csr_translator:av_readdata
	wire         atof_0_in_translator_avalon_anti_slave_0_waitrequest;                                               // atof_0:avalonmm_write_slave_waitrequest -> atof_0_in_translator:av_waitrequest
	wire  [31:0] atof_0_in_translator_avalon_anti_slave_0_writedata;                                                 // atof_0_in_translator:av_writedata -> atof_0:avalonmm_write_slave_writedata
	wire         atof_0_in_translator_avalon_anti_slave_0_write;                                                     // atof_0_in_translator:av_write -> atof_0:avalonmm_write_slave_write
	wire  [31:0] atof_0_in_csr_translator_avalon_anti_slave_0_writedata;                                             // atof_0_in_csr_translator:av_writedata -> atof_0:wrclk_control_slave_writedata
	wire   [2:0] atof_0_in_csr_translator_avalon_anti_slave_0_address;                                               // atof_0_in_csr_translator:av_address -> atof_0:wrclk_control_slave_address
	wire         atof_0_in_csr_translator_avalon_anti_slave_0_write;                                                 // atof_0_in_csr_translator:av_write -> atof_0:wrclk_control_slave_write
	wire         atof_0_in_csr_translator_avalon_anti_slave_0_read;                                                  // atof_0_in_csr_translator:av_read -> atof_0:wrclk_control_slave_read
	wire  [31:0] atof_0_in_csr_translator_avalon_anti_slave_0_readdata;                                              // atof_0:wrclk_control_slave_readdata -> atof_0_in_csr_translator:av_readdata
	wire         atof_0_out_translator_avalon_anti_slave_0_waitrequest;                                              // atof_0:avalonmm_read_slave_waitrequest -> atof_0_out_translator:av_waitrequest
	wire         atof_0_out_translator_avalon_anti_slave_0_read;                                                     // atof_0_out_translator:av_read -> atof_0:avalonmm_read_slave_read
	wire  [31:0] atof_0_out_translator_avalon_anti_slave_0_readdata;                                                 // atof_0:avalonmm_read_slave_readdata -> atof_0_out_translator:av_readdata
	wire  [31:0] ins_mem_5_s1_translator_avalon_anti_slave_0_writedata;                                              // ins_mem_5_s1_translator:av_writedata -> ins_mem_5:writedata
	wire   [9:0] ins_mem_5_s1_translator_avalon_anti_slave_0_address;                                                // ins_mem_5_s1_translator:av_address -> ins_mem_5:address
	wire         ins_mem_5_s1_translator_avalon_anti_slave_0_chipselect;                                             // ins_mem_5_s1_translator:av_chipselect -> ins_mem_5:chipselect
	wire         ins_mem_5_s1_translator_avalon_anti_slave_0_clken;                                                  // ins_mem_5_s1_translator:av_clken -> ins_mem_5:clken
	wire         ins_mem_5_s1_translator_avalon_anti_slave_0_write;                                                  // ins_mem_5_s1_translator:av_write -> ins_mem_5:write
	wire  [31:0] ins_mem_5_s1_translator_avalon_anti_slave_0_readdata;                                               // ins_mem_5:readdata -> ins_mem_5_s1_translator:av_readdata
	wire   [3:0] ins_mem_5_s1_translator_avalon_anti_slave_0_byteenable;                                             // ins_mem_5_s1_translator:av_byteenable -> ins_mem_5:byteenable
	wire  [31:0] cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_5_jtag_debug_module_translator:av_writedata -> cpu_5:jtag_debug_module_writedata
	wire   [8:0] cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_5_jtag_debug_module_translator:av_address -> cpu_5:jtag_debug_module_address
	wire         cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_5_jtag_debug_module_translator:av_chipselect -> cpu_5:jtag_debug_module_select
	wire         cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_5_jtag_debug_module_translator:av_write -> cpu_5:jtag_debug_module_write
	wire  [31:0] cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_5:jtag_debug_module_readdata -> cpu_5_jtag_debug_module_translator:av_readdata
	wire         cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_5_jtag_debug_module_translator:av_begintransfer -> cpu_5:jtag_debug_module_begintransfer
	wire         cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_5_jtag_debug_module_translator:av_debugaccess -> cpu_5:jtag_debug_module_debugaccess
	wire   [3:0] cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_5_jtag_debug_module_translator:av_byteenable -> cpu_5:jtag_debug_module_byteenable
	wire         etof_0_in_translator_avalon_anti_slave_0_waitrequest;                                               // etof_0:avalonmm_write_slave_waitrequest -> etof_0_in_translator:av_waitrequest
	wire  [31:0] etof_0_in_translator_avalon_anti_slave_0_writedata;                                                 // etof_0_in_translator:av_writedata -> etof_0:avalonmm_write_slave_writedata
	wire         etof_0_in_translator_avalon_anti_slave_0_write;                                                     // etof_0_in_translator:av_write -> etof_0:avalonmm_write_slave_write
	wire  [31:0] etof_0_in_csr_translator_avalon_anti_slave_0_writedata;                                             // etof_0_in_csr_translator:av_writedata -> etof_0:wrclk_control_slave_writedata
	wire   [2:0] etof_0_in_csr_translator_avalon_anti_slave_0_address;                                               // etof_0_in_csr_translator:av_address -> etof_0:wrclk_control_slave_address
	wire         etof_0_in_csr_translator_avalon_anti_slave_0_write;                                                 // etof_0_in_csr_translator:av_write -> etof_0:wrclk_control_slave_write
	wire         etof_0_in_csr_translator_avalon_anti_slave_0_read;                                                  // etof_0_in_csr_translator:av_read -> etof_0:wrclk_control_slave_read
	wire  [31:0] etof_0_in_csr_translator_avalon_anti_slave_0_readdata;                                              // etof_0:wrclk_control_slave_readdata -> etof_0_in_csr_translator:av_readdata
	wire         etof_0_out_translator_avalon_anti_slave_0_waitrequest;                                              // etof_0:avalonmm_read_slave_waitrequest -> etof_0_out_translator:av_waitrequest
	wire         etof_0_out_translator_avalon_anti_slave_0_read;                                                     // etof_0_out_translator:av_read -> etof_0:avalonmm_read_slave_read
	wire  [31:0] etof_0_out_translator_avalon_anti_slave_0_readdata;                                                 // etof_0:avalonmm_read_slave_readdata -> etof_0_out_translator:av_readdata
	wire  [31:0] data_mem_5_s1_translator_avalon_anti_slave_0_writedata;                                             // data_mem_5_s1_translator:av_writedata -> data_mem_5:writedata
	wire   [8:0] data_mem_5_s1_translator_avalon_anti_slave_0_address;                                               // data_mem_5_s1_translator:av_address -> data_mem_5:address
	wire         data_mem_5_s1_translator_avalon_anti_slave_0_chipselect;                                            // data_mem_5_s1_translator:av_chipselect -> data_mem_5:chipselect
	wire         data_mem_5_s1_translator_avalon_anti_slave_0_clken;                                                 // data_mem_5_s1_translator:av_clken -> data_mem_5:clken
	wire         data_mem_5_s1_translator_avalon_anti_slave_0_write;                                                 // data_mem_5_s1_translator:av_write -> data_mem_5:write
	wire  [31:0] data_mem_5_s1_translator_avalon_anti_slave_0_readdata;                                              // data_mem_5:readdata -> data_mem_5_s1_translator:av_readdata
	wire   [3:0] data_mem_5_s1_translator_avalon_anti_slave_0_byteenable;                                            // data_mem_5_s1_translator:av_byteenable -> data_mem_5:byteenable
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_5:av_waitrequest -> jtag_uart_5_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_5_avalon_jtag_slave_translator:av_writedata -> jtag_uart_5:av_writedata
	wire   [0:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_5_avalon_jtag_slave_translator:av_address -> jtag_uart_5:av_address
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_5_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_5:av_chipselect
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_5_avalon_jtag_slave_translator:av_write -> jtag_uart_5:av_write_n
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_5_avalon_jtag_slave_translator:av_read -> jtag_uart_5:av_read_n
	wire  [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_5:av_readdata -> jtag_uart_5_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_5_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_5_s1_translator:av_writedata -> timer_5:writedata
	wire   [2:0] timer_5_s1_translator_avalon_anti_slave_0_address;                                                  // timer_5_s1_translator:av_address -> timer_5:address
	wire         timer_5_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_5_s1_translator:av_chipselect -> timer_5:chipselect
	wire         timer_5_s1_translator_avalon_anti_slave_0_write;                                                    // timer_5_s1_translator:av_write -> timer_5:write_n
	wire  [15:0] timer_5_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_5:readdata -> timer_5_s1_translator:av_readdata
	wire  [15:0] high_scale_timer_5_s1_translator_avalon_anti_slave_0_writedata;                                     // high_scale_timer_5_s1_translator:av_writedata -> high_scale_timer_5:writedata
	wire   [2:0] high_scale_timer_5_s1_translator_avalon_anti_slave_0_address;                                       // high_scale_timer_5_s1_translator:av_address -> high_scale_timer_5:address
	wire         high_scale_timer_5_s1_translator_avalon_anti_slave_0_chipselect;                                    // high_scale_timer_5_s1_translator:av_chipselect -> high_scale_timer_5:chipselect
	wire         high_scale_timer_5_s1_translator_avalon_anti_slave_0_write;                                         // high_scale_timer_5_s1_translator:av_write -> high_scale_timer_5:write_n
	wire  [15:0] high_scale_timer_5_s1_translator_avalon_anti_slave_0_readdata;                                      // high_scale_timer_5:readdata -> high_scale_timer_5_s1_translator:av_readdata
	wire  [31:0] data_mem_0_s1_translator_avalon_anti_slave_0_writedata;                                             // data_mem_0_s1_translator:av_writedata -> data_mem_0:writedata
	wire   [8:0] data_mem_0_s1_translator_avalon_anti_slave_0_address;                                               // data_mem_0_s1_translator:av_address -> data_mem_0:address
	wire         data_mem_0_s1_translator_avalon_anti_slave_0_chipselect;                                            // data_mem_0_s1_translator:av_chipselect -> data_mem_0:chipselect
	wire         data_mem_0_s1_translator_avalon_anti_slave_0_clken;                                                 // data_mem_0_s1_translator:av_clken -> data_mem_0:clken
	wire         data_mem_0_s1_translator_avalon_anti_slave_0_write;                                                 // data_mem_0_s1_translator:av_write -> data_mem_0:write
	wire  [31:0] data_mem_0_s1_translator_avalon_anti_slave_0_readdata;                                              // data_mem_0:readdata -> data_mem_0_s1_translator:av_readdata
	wire   [3:0] data_mem_0_s1_translator_avalon_anti_slave_0_byteenable;                                            // data_mem_0_s1_translator:av_byteenable -> data_mem_0:byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                  // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                    // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire  [15:0] high_scale_timer_0_s1_translator_avalon_anti_slave_0_writedata;                                     // high_scale_timer_0_s1_translator:av_writedata -> high_scale_timer_0:writedata
	wire   [2:0] high_scale_timer_0_s1_translator_avalon_anti_slave_0_address;                                       // high_scale_timer_0_s1_translator:av_address -> high_scale_timer_0:address
	wire         high_scale_timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                    // high_scale_timer_0_s1_translator:av_chipselect -> high_scale_timer_0:chipselect
	wire         high_scale_timer_0_s1_translator_avalon_anti_slave_0_write;                                         // high_scale_timer_0_s1_translator:av_write -> high_scale_timer_0:write_n
	wire  [15:0] high_scale_timer_0_s1_translator_avalon_anti_slave_0_readdata;                                      // high_scale_timer_0:readdata -> high_scale_timer_0_s1_translator:av_readdata
	wire  [31:0] ins_mem_4_s1_translator_avalon_anti_slave_0_writedata;                                              // ins_mem_4_s1_translator:av_writedata -> ins_mem_4:writedata
	wire   [9:0] ins_mem_4_s1_translator_avalon_anti_slave_0_address;                                                // ins_mem_4_s1_translator:av_address -> ins_mem_4:address
	wire         ins_mem_4_s1_translator_avalon_anti_slave_0_chipselect;                                             // ins_mem_4_s1_translator:av_chipselect -> ins_mem_4:chipselect
	wire         ins_mem_4_s1_translator_avalon_anti_slave_0_clken;                                                  // ins_mem_4_s1_translator:av_clken -> ins_mem_4:clken
	wire         ins_mem_4_s1_translator_avalon_anti_slave_0_write;                                                  // ins_mem_4_s1_translator:av_write -> ins_mem_4:write
	wire  [31:0] ins_mem_4_s1_translator_avalon_anti_slave_0_readdata;                                               // ins_mem_4:readdata -> ins_mem_4_s1_translator:av_readdata
	wire   [3:0] ins_mem_4_s1_translator_avalon_anti_slave_0_byteenable;                                             // ins_mem_4_s1_translator:av_byteenable -> ins_mem_4:byteenable
	wire  [31:0] cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_4_jtag_debug_module_translator:av_writedata -> cpu_4:jtag_debug_module_writedata
	wire   [8:0] cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_4_jtag_debug_module_translator:av_address -> cpu_4:jtag_debug_module_address
	wire         cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_4_jtag_debug_module_translator:av_chipselect -> cpu_4:jtag_debug_module_select
	wire         cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_4_jtag_debug_module_translator:av_write -> cpu_4:jtag_debug_module_write
	wire  [31:0] cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_4:jtag_debug_module_readdata -> cpu_4_jtag_debug_module_translator:av_readdata
	wire         cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_4_jtag_debug_module_translator:av_begintransfer -> cpu_4:jtag_debug_module_begintransfer
	wire         cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_4_jtag_debug_module_translator:av_debugaccess -> cpu_4:jtag_debug_module_debugaccess
	wire   [3:0] cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_4_jtag_debug_module_translator:av_byteenable -> cpu_4:jtag_debug_module_byteenable
	wire         dtoe_0_in_translator_avalon_anti_slave_0_waitrequest;                                               // dtoe_0:avalonmm_write_slave_waitrequest -> dtoe_0_in_translator:av_waitrequest
	wire  [31:0] dtoe_0_in_translator_avalon_anti_slave_0_writedata;                                                 // dtoe_0_in_translator:av_writedata -> dtoe_0:avalonmm_write_slave_writedata
	wire         dtoe_0_in_translator_avalon_anti_slave_0_write;                                                     // dtoe_0_in_translator:av_write -> dtoe_0:avalonmm_write_slave_write
	wire  [31:0] dtoe_0_in_csr_translator_avalon_anti_slave_0_writedata;                                             // dtoe_0_in_csr_translator:av_writedata -> dtoe_0:wrclk_control_slave_writedata
	wire   [2:0] dtoe_0_in_csr_translator_avalon_anti_slave_0_address;                                               // dtoe_0_in_csr_translator:av_address -> dtoe_0:wrclk_control_slave_address
	wire         dtoe_0_in_csr_translator_avalon_anti_slave_0_write;                                                 // dtoe_0_in_csr_translator:av_write -> dtoe_0:wrclk_control_slave_write
	wire         dtoe_0_in_csr_translator_avalon_anti_slave_0_read;                                                  // dtoe_0_in_csr_translator:av_read -> dtoe_0:wrclk_control_slave_read
	wire  [31:0] dtoe_0_in_csr_translator_avalon_anti_slave_0_readdata;                                              // dtoe_0:wrclk_control_slave_readdata -> dtoe_0_in_csr_translator:av_readdata
	wire         dtoe_0_out_translator_avalon_anti_slave_0_waitrequest;                                              // dtoe_0:avalonmm_read_slave_waitrequest -> dtoe_0_out_translator:av_waitrequest
	wire         dtoe_0_out_translator_avalon_anti_slave_0_read;                                                     // dtoe_0_out_translator:av_read -> dtoe_0:avalonmm_read_slave_read
	wire  [31:0] dtoe_0_out_translator_avalon_anti_slave_0_readdata;                                                 // dtoe_0:avalonmm_read_slave_readdata -> dtoe_0_out_translator:av_readdata
	wire  [31:0] data_mem_4_s1_translator_avalon_anti_slave_0_writedata;                                             // data_mem_4_s1_translator:av_writedata -> data_mem_4:writedata
	wire   [8:0] data_mem_4_s1_translator_avalon_anti_slave_0_address;                                               // data_mem_4_s1_translator:av_address -> data_mem_4:address
	wire         data_mem_4_s1_translator_avalon_anti_slave_0_chipselect;                                            // data_mem_4_s1_translator:av_chipselect -> data_mem_4:chipselect
	wire         data_mem_4_s1_translator_avalon_anti_slave_0_clken;                                                 // data_mem_4_s1_translator:av_clken -> data_mem_4:clken
	wire         data_mem_4_s1_translator_avalon_anti_slave_0_write;                                                 // data_mem_4_s1_translator:av_write -> data_mem_4:write
	wire  [31:0] data_mem_4_s1_translator_avalon_anti_slave_0_readdata;                                              // data_mem_4:readdata -> data_mem_4_s1_translator:av_readdata
	wire   [3:0] data_mem_4_s1_translator_avalon_anti_slave_0_byteenable;                                            // data_mem_4_s1_translator:av_byteenable -> data_mem_4:byteenable
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_4:av_waitrequest -> jtag_uart_4_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_4_avalon_jtag_slave_translator:av_writedata -> jtag_uart_4:av_writedata
	wire   [0:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_4_avalon_jtag_slave_translator:av_address -> jtag_uart_4:av_address
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_4_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_4:av_chipselect
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_4_avalon_jtag_slave_translator:av_write -> jtag_uart_4:av_write_n
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_4_avalon_jtag_slave_translator:av_read -> jtag_uart_4:av_read_n
	wire  [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_4:av_readdata -> jtag_uart_4_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_4_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_4_s1_translator:av_writedata -> timer_4:writedata
	wire   [2:0] timer_4_s1_translator_avalon_anti_slave_0_address;                                                  // timer_4_s1_translator:av_address -> timer_4:address
	wire         timer_4_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_4_s1_translator:av_chipselect -> timer_4:chipselect
	wire         timer_4_s1_translator_avalon_anti_slave_0_write;                                                    // timer_4_s1_translator:av_write -> timer_4:write_n
	wire  [15:0] timer_4_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_4:readdata -> timer_4_s1_translator:av_readdata
	wire  [15:0] high_scale_timer_4_s1_translator_avalon_anti_slave_0_writedata;                                     // high_scale_timer_4_s1_translator:av_writedata -> high_scale_timer_4:writedata
	wire   [2:0] high_scale_timer_4_s1_translator_avalon_anti_slave_0_address;                                       // high_scale_timer_4_s1_translator:av_address -> high_scale_timer_4:address
	wire         high_scale_timer_4_s1_translator_avalon_anti_slave_0_chipselect;                                    // high_scale_timer_4_s1_translator:av_chipselect -> high_scale_timer_4:chipselect
	wire         high_scale_timer_4_s1_translator_avalon_anti_slave_0_write;                                         // high_scale_timer_4_s1_translator:av_write -> high_scale_timer_4:write_n
	wire  [15:0] high_scale_timer_4_s1_translator_avalon_anti_slave_0_readdata;                                      // high_scale_timer_4:readdata -> high_scale_timer_4_s1_translator:av_readdata
	wire  [31:0] ins_mem_3_s1_translator_avalon_anti_slave_0_writedata;                                              // ins_mem_3_s1_translator:av_writedata -> ins_mem_3:writedata
	wire   [9:0] ins_mem_3_s1_translator_avalon_anti_slave_0_address;                                                // ins_mem_3_s1_translator:av_address -> ins_mem_3:address
	wire         ins_mem_3_s1_translator_avalon_anti_slave_0_chipselect;                                             // ins_mem_3_s1_translator:av_chipselect -> ins_mem_3:chipselect
	wire         ins_mem_3_s1_translator_avalon_anti_slave_0_clken;                                                  // ins_mem_3_s1_translator:av_clken -> ins_mem_3:clken
	wire         ins_mem_3_s1_translator_avalon_anti_slave_0_write;                                                  // ins_mem_3_s1_translator:av_write -> ins_mem_3:write
	wire  [31:0] ins_mem_3_s1_translator_avalon_anti_slave_0_readdata;                                               // ins_mem_3:readdata -> ins_mem_3_s1_translator:av_readdata
	wire   [3:0] ins_mem_3_s1_translator_avalon_anti_slave_0_byteenable;                                             // ins_mem_3_s1_translator:av_byteenable -> ins_mem_3:byteenable
	wire  [31:0] cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_3_jtag_debug_module_translator:av_writedata -> cpu_3:jtag_debug_module_writedata
	wire   [8:0] cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_3_jtag_debug_module_translator:av_address -> cpu_3:jtag_debug_module_address
	wire         cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_3_jtag_debug_module_translator:av_chipselect -> cpu_3:jtag_debug_module_select
	wire         cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_3_jtag_debug_module_translator:av_write -> cpu_3:jtag_debug_module_write
	wire  [31:0] cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_3:jtag_debug_module_readdata -> cpu_3_jtag_debug_module_translator:av_readdata
	wire         cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_3_jtag_debug_module_translator:av_begintransfer -> cpu_3:jtag_debug_module_begintransfer
	wire         cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_3_jtag_debug_module_translator:av_debugaccess -> cpu_3:jtag_debug_module_debugaccess
	wire   [3:0] cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_3_jtag_debug_module_translator:av_byteenable -> cpu_3:jtag_debug_module_byteenable
	wire         ctod_0_in_translator_avalon_anti_slave_0_waitrequest;                                               // ctod_0:avalonmm_write_slave_waitrequest -> ctod_0_in_translator:av_waitrequest
	wire  [31:0] ctod_0_in_translator_avalon_anti_slave_0_writedata;                                                 // ctod_0_in_translator:av_writedata -> ctod_0:avalonmm_write_slave_writedata
	wire         ctod_0_in_translator_avalon_anti_slave_0_write;                                                     // ctod_0_in_translator:av_write -> ctod_0:avalonmm_write_slave_write
	wire  [31:0] ctod_0_in_csr_translator_avalon_anti_slave_0_writedata;                                             // ctod_0_in_csr_translator:av_writedata -> ctod_0:wrclk_control_slave_writedata
	wire   [2:0] ctod_0_in_csr_translator_avalon_anti_slave_0_address;                                               // ctod_0_in_csr_translator:av_address -> ctod_0:wrclk_control_slave_address
	wire         ctod_0_in_csr_translator_avalon_anti_slave_0_write;                                                 // ctod_0_in_csr_translator:av_write -> ctod_0:wrclk_control_slave_write
	wire         ctod_0_in_csr_translator_avalon_anti_slave_0_read;                                                  // ctod_0_in_csr_translator:av_read -> ctod_0:wrclk_control_slave_read
	wire  [31:0] ctod_0_in_csr_translator_avalon_anti_slave_0_readdata;                                              // ctod_0:wrclk_control_slave_readdata -> ctod_0_in_csr_translator:av_readdata
	wire         ctod_0_out_translator_avalon_anti_slave_0_waitrequest;                                              // ctod_0:avalonmm_read_slave_waitrequest -> ctod_0_out_translator:av_waitrequest
	wire         ctod_0_out_translator_avalon_anti_slave_0_read;                                                     // ctod_0_out_translator:av_read -> ctod_0:avalonmm_read_slave_read
	wire  [31:0] ctod_0_out_translator_avalon_anti_slave_0_readdata;                                                 // ctod_0:avalonmm_read_slave_readdata -> ctod_0_out_translator:av_readdata
	wire  [31:0] data_mem_3_s1_translator_avalon_anti_slave_0_writedata;                                             // data_mem_3_s1_translator:av_writedata -> data_mem_3:writedata
	wire   [8:0] data_mem_3_s1_translator_avalon_anti_slave_0_address;                                               // data_mem_3_s1_translator:av_address -> data_mem_3:address
	wire         data_mem_3_s1_translator_avalon_anti_slave_0_chipselect;                                            // data_mem_3_s1_translator:av_chipselect -> data_mem_3:chipselect
	wire         data_mem_3_s1_translator_avalon_anti_slave_0_clken;                                                 // data_mem_3_s1_translator:av_clken -> data_mem_3:clken
	wire         data_mem_3_s1_translator_avalon_anti_slave_0_write;                                                 // data_mem_3_s1_translator:av_write -> data_mem_3:write
	wire  [31:0] data_mem_3_s1_translator_avalon_anti_slave_0_readdata;                                              // data_mem_3:readdata -> data_mem_3_s1_translator:av_readdata
	wire   [3:0] data_mem_3_s1_translator_avalon_anti_slave_0_byteenable;                                            // data_mem_3_s1_translator:av_byteenable -> data_mem_3:byteenable
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_3:av_waitrequest -> jtag_uart_3_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_3_avalon_jtag_slave_translator:av_writedata -> jtag_uart_3:av_writedata
	wire   [0:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_3_avalon_jtag_slave_translator:av_address -> jtag_uart_3:av_address
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_3_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_3:av_chipselect
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_3_avalon_jtag_slave_translator:av_write -> jtag_uart_3:av_write_n
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_3_avalon_jtag_slave_translator:av_read -> jtag_uart_3:av_read_n
	wire  [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_3:av_readdata -> jtag_uart_3_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_3_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_3_s1_translator:av_writedata -> timer_3:writedata
	wire   [2:0] timer_3_s1_translator_avalon_anti_slave_0_address;                                                  // timer_3_s1_translator:av_address -> timer_3:address
	wire         timer_3_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_3_s1_translator:av_chipselect -> timer_3:chipselect
	wire         timer_3_s1_translator_avalon_anti_slave_0_write;                                                    // timer_3_s1_translator:av_write -> timer_3:write_n
	wire  [15:0] timer_3_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_3:readdata -> timer_3_s1_translator:av_readdata
	wire  [15:0] high_scale_timer_3_s1_translator_avalon_anti_slave_0_writedata;                                     // high_scale_timer_3_s1_translator:av_writedata -> high_scale_timer_3:writedata
	wire   [2:0] high_scale_timer_3_s1_translator_avalon_anti_slave_0_address;                                       // high_scale_timer_3_s1_translator:av_address -> high_scale_timer_3:address
	wire         high_scale_timer_3_s1_translator_avalon_anti_slave_0_chipselect;                                    // high_scale_timer_3_s1_translator:av_chipselect -> high_scale_timer_3:chipselect
	wire         high_scale_timer_3_s1_translator_avalon_anti_slave_0_write;                                         // high_scale_timer_3_s1_translator:av_write -> high_scale_timer_3:write_n
	wire  [15:0] high_scale_timer_3_s1_translator_avalon_anti_slave_0_readdata;                                      // high_scale_timer_3:readdata -> high_scale_timer_3_s1_translator:av_readdata
	wire  [31:0] data_mem_2_s1_translator_avalon_anti_slave_0_writedata;                                             // data_mem_2_s1_translator:av_writedata -> data_mem_2:writedata
	wire   [8:0] data_mem_2_s1_translator_avalon_anti_slave_0_address;                                               // data_mem_2_s1_translator:av_address -> data_mem_2:address
	wire         data_mem_2_s1_translator_avalon_anti_slave_0_chipselect;                                            // data_mem_2_s1_translator:av_chipselect -> data_mem_2:chipselect
	wire         data_mem_2_s1_translator_avalon_anti_slave_0_clken;                                                 // data_mem_2_s1_translator:av_clken -> data_mem_2:clken
	wire         data_mem_2_s1_translator_avalon_anti_slave_0_write;                                                 // data_mem_2_s1_translator:av_write -> data_mem_2:write
	wire  [31:0] data_mem_2_s1_translator_avalon_anti_slave_0_readdata;                                              // data_mem_2:readdata -> data_mem_2_s1_translator:av_readdata
	wire   [3:0] data_mem_2_s1_translator_avalon_anti_slave_0_byteenable;                                            // data_mem_2_s1_translator:av_byteenable -> data_mem_2:byteenable
	wire  [31:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_2_jtag_debug_module_translator:av_writedata -> cpu_2:jtag_debug_module_writedata
	wire   [8:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_2_jtag_debug_module_translator:av_address -> cpu_2:jtag_debug_module_address
	wire         cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_2_jtag_debug_module_translator:av_chipselect -> cpu_2:jtag_debug_module_select
	wire         cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_2_jtag_debug_module_translator:av_write -> cpu_2:jtag_debug_module_write
	wire  [31:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_2:jtag_debug_module_readdata -> cpu_2_jtag_debug_module_translator:av_readdata
	wire         cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_2_jtag_debug_module_translator:av_begintransfer -> cpu_2:jtag_debug_module_begintransfer
	wire         cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_2_jtag_debug_module_translator:av_debugaccess -> cpu_2:jtag_debug_module_debugaccess
	wire   [3:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_2_jtag_debug_module_translator:av_byteenable -> cpu_2:jtag_debug_module_byteenable
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_2:av_waitrequest -> jtag_uart_2_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_2_avalon_jtag_slave_translator:av_writedata -> jtag_uart_2:av_writedata
	wire   [0:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_2_avalon_jtag_slave_translator:av_address -> jtag_uart_2:av_address
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_2_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_2:av_chipselect
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_2_avalon_jtag_slave_translator:av_write -> jtag_uart_2:av_write_n
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_2_avalon_jtag_slave_translator:av_read -> jtag_uart_2:av_read_n
	wire  [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_2:av_readdata -> jtag_uart_2_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_2_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_2_s1_translator:av_writedata -> timer_2:writedata
	wire   [2:0] timer_2_s1_translator_avalon_anti_slave_0_address;                                                  // timer_2_s1_translator:av_address -> timer_2:address
	wire         timer_2_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_2_s1_translator:av_chipselect -> timer_2:chipselect
	wire         timer_2_s1_translator_avalon_anti_slave_0_write;                                                    // timer_2_s1_translator:av_write -> timer_2:write_n
	wire  [15:0] timer_2_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_2:readdata -> timer_2_s1_translator:av_readdata
	wire  [15:0] high_scale_timer_2_s1_translator_avalon_anti_slave_0_writedata;                                     // high_scale_timer_2_s1_translator:av_writedata -> high_scale_timer_2:writedata
	wire   [2:0] high_scale_timer_2_s1_translator_avalon_anti_slave_0_address;                                       // high_scale_timer_2_s1_translator:av_address -> high_scale_timer_2:address
	wire         high_scale_timer_2_s1_translator_avalon_anti_slave_0_chipselect;                                    // high_scale_timer_2_s1_translator:av_chipselect -> high_scale_timer_2:chipselect
	wire         high_scale_timer_2_s1_translator_avalon_anti_slave_0_write;                                         // high_scale_timer_2_s1_translator:av_write -> high_scale_timer_2:write_n
	wire  [15:0] high_scale_timer_2_s1_translator_avalon_anti_slave_0_readdata;                                      // high_scale_timer_2:readdata -> high_scale_timer_2_s1_translator:av_readdata
	wire         btoc_0_in_translator_avalon_anti_slave_0_waitrequest;                                               // btoc_0:avalonmm_write_slave_waitrequest -> btoc_0_in_translator:av_waitrequest
	wire  [31:0] btoc_0_in_translator_avalon_anti_slave_0_writedata;                                                 // btoc_0_in_translator:av_writedata -> btoc_0:avalonmm_write_slave_writedata
	wire         btoc_0_in_translator_avalon_anti_slave_0_write;                                                     // btoc_0_in_translator:av_write -> btoc_0:avalonmm_write_slave_write
	wire         btoc_0_out_translator_avalon_anti_slave_0_waitrequest;                                              // btoc_0:avalonmm_read_slave_waitrequest -> btoc_0_out_translator:av_waitrequest
	wire         btoc_0_out_translator_avalon_anti_slave_0_read;                                                     // btoc_0_out_translator:av_read -> btoc_0:avalonmm_read_slave_read
	wire  [31:0] btoc_0_out_translator_avalon_anti_slave_0_readdata;                                                 // btoc_0:avalonmm_read_slave_readdata -> btoc_0_out_translator:av_readdata
	wire  [31:0] btoc_0_in_csr_translator_avalon_anti_slave_0_writedata;                                             // btoc_0_in_csr_translator:av_writedata -> btoc_0:wrclk_control_slave_writedata
	wire   [2:0] btoc_0_in_csr_translator_avalon_anti_slave_0_address;                                               // btoc_0_in_csr_translator:av_address -> btoc_0:wrclk_control_slave_address
	wire         btoc_0_in_csr_translator_avalon_anti_slave_0_write;                                                 // btoc_0_in_csr_translator:av_write -> btoc_0:wrclk_control_slave_write
	wire         btoc_0_in_csr_translator_avalon_anti_slave_0_read;                                                  // btoc_0_in_csr_translator:av_read -> btoc_0:wrclk_control_slave_read
	wire  [31:0] btoc_0_in_csr_translator_avalon_anti_slave_0_readdata;                                              // btoc_0:wrclk_control_slave_readdata -> btoc_0_in_csr_translator:av_readdata
	wire  [31:0] ins_mem_2_s1_translator_avalon_anti_slave_0_writedata;                                              // ins_mem_2_s1_translator:av_writedata -> ins_mem_2:writedata
	wire   [9:0] ins_mem_2_s1_translator_avalon_anti_slave_0_address;                                                // ins_mem_2_s1_translator:av_address -> ins_mem_2:address
	wire         ins_mem_2_s1_translator_avalon_anti_slave_0_chipselect;                                             // ins_mem_2_s1_translator:av_chipselect -> ins_mem_2:chipselect
	wire         ins_mem_2_s1_translator_avalon_anti_slave_0_clken;                                                  // ins_mem_2_s1_translator:av_clken -> ins_mem_2:clken
	wire         ins_mem_2_s1_translator_avalon_anti_slave_0_write;                                                  // ins_mem_2_s1_translator:av_write -> ins_mem_2:write
	wire  [31:0] ins_mem_2_s1_translator_avalon_anti_slave_0_readdata;                                               // ins_mem_2:readdata -> ins_mem_2_s1_translator:av_readdata
	wire   [3:0] ins_mem_2_s1_translator_avalon_anti_slave_0_byteenable;                                             // ins_mem_2_s1_translator:av_byteenable -> ins_mem_2:byteenable
	wire  [31:0] ins_mem_1_s1_translator_avalon_anti_slave_0_writedata;                                              // ins_mem_1_s1_translator:av_writedata -> ins_mem_1:writedata
	wire   [9:0] ins_mem_1_s1_translator_avalon_anti_slave_0_address;                                                // ins_mem_1_s1_translator:av_address -> ins_mem_1:address
	wire         ins_mem_1_s1_translator_avalon_anti_slave_0_chipselect;                                             // ins_mem_1_s1_translator:av_chipselect -> ins_mem_1:chipselect
	wire         ins_mem_1_s1_translator_avalon_anti_slave_0_clken;                                                  // ins_mem_1_s1_translator:av_clken -> ins_mem_1:clken
	wire         ins_mem_1_s1_translator_avalon_anti_slave_0_write;                                                  // ins_mem_1_s1_translator:av_write -> ins_mem_1:write
	wire  [31:0] ins_mem_1_s1_translator_avalon_anti_slave_0_readdata;                                               // ins_mem_1:readdata -> ins_mem_1_s1_translator:av_readdata
	wire   [3:0] ins_mem_1_s1_translator_avalon_anti_slave_0_byteenable;                                             // ins_mem_1_s1_translator:av_byteenable -> ins_mem_1:byteenable
	wire  [31:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_1_jtag_debug_module_translator:av_writedata -> cpu_1:jtag_debug_module_writedata
	wire   [8:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_1_jtag_debug_module_translator:av_address -> cpu_1:jtag_debug_module_address
	wire         cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                  // cpu_1_jtag_debug_module_translator:av_chipselect -> cpu_1:jtag_debug_module_select
	wire         cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_1_jtag_debug_module_translator:av_write -> cpu_1:jtag_debug_module_write
	wire  [31:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu_1:jtag_debug_module_readdata -> cpu_1_jtag_debug_module_translator:av_readdata
	wire         cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                               // cpu_1_jtag_debug_module_translator:av_begintransfer -> cpu_1:jtag_debug_module_begintransfer
	wire         cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_1_jtag_debug_module_translator:av_debugaccess -> cpu_1:jtag_debug_module_debugaccess
	wire   [3:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_1_jtag_debug_module_translator:av_byteenable -> cpu_1:jtag_debug_module_byteenable
	wire  [31:0] data_mem_1_s1_translator_avalon_anti_slave_0_writedata;                                             // data_mem_1_s1_translator:av_writedata -> data_mem_1:writedata
	wire   [8:0] data_mem_1_s1_translator_avalon_anti_slave_0_address;                                               // data_mem_1_s1_translator:av_address -> data_mem_1:address
	wire         data_mem_1_s1_translator_avalon_anti_slave_0_chipselect;                                            // data_mem_1_s1_translator:av_chipselect -> data_mem_1:chipselect
	wire         data_mem_1_s1_translator_avalon_anti_slave_0_clken;                                                 // data_mem_1_s1_translator:av_clken -> data_mem_1:clken
	wire         data_mem_1_s1_translator_avalon_anti_slave_0_write;                                                 // data_mem_1_s1_translator:av_write -> data_mem_1:write
	wire  [31:0] data_mem_1_s1_translator_avalon_anti_slave_0_readdata;                                              // data_mem_1:readdata -> data_mem_1_s1_translator:av_readdata
	wire   [3:0] data_mem_1_s1_translator_avalon_anti_slave_0_byteenable;                                            // data_mem_1_s1_translator:av_byteenable -> data_mem_1:byteenable
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_1:av_waitrequest -> jtag_uart_1_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_1_avalon_jtag_slave_translator:av_writedata -> jtag_uart_1:av_writedata
	wire   [0:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_1_avalon_jtag_slave_translator:av_address -> jtag_uart_1:av_address
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_1_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_1:av_chipselect
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_1_avalon_jtag_slave_translator:av_write -> jtag_uart_1:av_write_n
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_1_avalon_jtag_slave_translator:av_read -> jtag_uart_1:av_read_n
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_1:av_readdata -> jtag_uart_1_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_1_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_1_s1_translator:av_writedata -> timer_1:writedata
	wire   [2:0] timer_1_s1_translator_avalon_anti_slave_0_address;                                                  // timer_1_s1_translator:av_address -> timer_1:address
	wire         timer_1_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	wire         timer_1_s1_translator_avalon_anti_slave_0_write;                                                    // timer_1_s1_translator:av_write -> timer_1:write_n
	wire  [15:0] timer_1_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_1:readdata -> timer_1_s1_translator:av_readdata
	wire  [15:0] high_scale_timer_1_s1_translator_avalon_anti_slave_0_writedata;                                     // high_scale_timer_1_s1_translator:av_writedata -> high_scale_timer_1:writedata
	wire   [2:0] high_scale_timer_1_s1_translator_avalon_anti_slave_0_address;                                       // high_scale_timer_1_s1_translator:av_address -> high_scale_timer_1:address
	wire         high_scale_timer_1_s1_translator_avalon_anti_slave_0_chipselect;                                    // high_scale_timer_1_s1_translator:av_chipselect -> high_scale_timer_1:chipselect
	wire         high_scale_timer_1_s1_translator_avalon_anti_slave_0_write;                                         // high_scale_timer_1_s1_translator:av_write -> high_scale_timer_1:write_n
	wire  [15:0] high_scale_timer_1_s1_translator_avalon_anti_slave_0_readdata;                                      // high_scale_timer_1:readdata -> high_scale_timer_1_s1_translator:av_readdata
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_0_instruction_master_translator:uav_burstcount -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_0_instruction_master_translator:uav_writedata -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_0_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_0_instruction_master_translator:uav_address -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_0_instruction_master_translator:uav_lock -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_0_instruction_master_translator:uav_write -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_0_instruction_master_translator:uav_read -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_instruction_master_translator:uav_readdata
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_0_instruction_master_translator:uav_debugaccess -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_0_instruction_master_translator:uav_byteenable -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_instruction_master_translator:uav_readdatavalid
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_5_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_5_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_5_instruction_master_translator:uav_burstcount -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_5_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_5_instruction_master_translator:uav_writedata -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_5_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_5_instruction_master_translator:uav_address -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_5_instruction_master_translator:uav_lock -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_5_instruction_master_translator:uav_write -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_5_instruction_master_translator:uav_read -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_5_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_5_instruction_master_translator:uav_readdata
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_5_instruction_master_translator:uav_debugaccess -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_5_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_5_instruction_master_translator:uav_byteenable -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_5_instruction_master_translator:uav_readdatavalid
	wire         cpu_5_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_5_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_5_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_5_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_5_data_master_translator:uav_burstcount -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_5_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_5_data_master_translator:uav_writedata -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_5_data_master_translator_avalon_universal_master_0_address;                                     // cpu_5_data_master_translator:uav_address -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_5_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_5_data_master_translator:uav_lock -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_5_data_master_translator_avalon_universal_master_0_write;                                       // cpu_5_data_master_translator:uav_write -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_5_data_master_translator_avalon_universal_master_0_read;                                        // cpu_5_data_master_translator:uav_read -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_5_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_5_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_5_data_master_translator:uav_readdata
	wire         cpu_5_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_5_data_master_translator:uav_debugaccess -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_5_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_5_data_master_translator:uav_byteenable -> cpu_5_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_5_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_5_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_5_data_master_translator:uav_readdatavalid
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_4_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_4_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_4_instruction_master_translator:uav_burstcount -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_4_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_4_instruction_master_translator:uav_writedata -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_4_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_4_instruction_master_translator:uav_address -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_4_instruction_master_translator:uav_lock -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_4_instruction_master_translator:uav_write -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_4_instruction_master_translator:uav_read -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_4_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_4_instruction_master_translator:uav_readdata
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_4_instruction_master_translator:uav_debugaccess -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_4_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_4_instruction_master_translator:uav_byteenable -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_4_instruction_master_translator:uav_readdatavalid
	wire         cpu_4_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_4_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_4_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_4_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_4_data_master_translator:uav_burstcount -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_4_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_4_data_master_translator:uav_writedata -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_4_data_master_translator_avalon_universal_master_0_address;                                     // cpu_4_data_master_translator:uav_address -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_4_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_4_data_master_translator:uav_lock -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_4_data_master_translator_avalon_universal_master_0_write;                                       // cpu_4_data_master_translator:uav_write -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_4_data_master_translator_avalon_universal_master_0_read;                                        // cpu_4_data_master_translator:uav_read -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_4_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_4_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_4_data_master_translator:uav_readdata
	wire         cpu_4_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_4_data_master_translator:uav_debugaccess -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_4_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_4_data_master_translator:uav_byteenable -> cpu_4_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_4_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_4_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_4_data_master_translator:uav_readdatavalid
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_3_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_3_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_3_instruction_master_translator:uav_burstcount -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_3_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_3_instruction_master_translator:uav_writedata -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_3_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_3_instruction_master_translator:uav_address -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_3_instruction_master_translator:uav_lock -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_3_instruction_master_translator:uav_write -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_3_instruction_master_translator:uav_read -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_3_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_3_instruction_master_translator:uav_readdata
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_3_instruction_master_translator:uav_debugaccess -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_3_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_3_instruction_master_translator:uav_byteenable -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_3_instruction_master_translator:uav_readdatavalid
	wire         cpu_3_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_3_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_3_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_3_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_3_data_master_translator:uav_burstcount -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_3_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_3_data_master_translator:uav_writedata -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_3_data_master_translator_avalon_universal_master_0_address;                                     // cpu_3_data_master_translator:uav_address -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_3_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_3_data_master_translator:uav_lock -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_3_data_master_translator_avalon_universal_master_0_write;                                       // cpu_3_data_master_translator:uav_write -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_3_data_master_translator_avalon_universal_master_0_read;                                        // cpu_3_data_master_translator:uav_read -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_3_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_3_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_3_data_master_translator:uav_readdata
	wire         cpu_3_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_3_data_master_translator:uav_debugaccess -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_3_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_3_data_master_translator:uav_byteenable -> cpu_3_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_3_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_3_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_3_data_master_translator:uav_readdatavalid
	wire         cpu_2_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_2_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_2_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_2_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_2_data_master_translator:uav_burstcount -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_2_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_2_data_master_translator:uav_writedata -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_2_data_master_translator_avalon_universal_master_0_address;                                     // cpu_2_data_master_translator:uav_address -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_2_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_2_data_master_translator:uav_lock -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_2_data_master_translator_avalon_universal_master_0_write;                                       // cpu_2_data_master_translator:uav_write -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_2_data_master_translator_avalon_universal_master_0_read;                                        // cpu_2_data_master_translator:uav_read -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_2_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_2_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_2_data_master_translator:uav_readdata
	wire         cpu_2_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_2_data_master_translator:uav_debugaccess -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_2_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_2_data_master_translator:uav_byteenable -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_2_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_2_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_2_data_master_translator:uav_readdatavalid
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_2_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_2_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_2_instruction_master_translator:uav_burstcount -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_2_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_2_instruction_master_translator:uav_writedata -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_2_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_2_instruction_master_translator:uav_address -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_2_instruction_master_translator:uav_lock -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_2_instruction_master_translator:uav_write -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_2_instruction_master_translator:uav_read -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_2_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_2_instruction_master_translator:uav_readdata
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_2_instruction_master_translator:uav_debugaccess -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_2_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_2_instruction_master_translator:uav_byteenable -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_2_instruction_master_translator:uav_readdatavalid
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_1_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_1_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_1_instruction_master_translator:uav_burstcount -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_1_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_1_instruction_master_translator:uav_writedata -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_1_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_1_instruction_master_translator:uav_address -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_1_instruction_master_translator:uav_lock -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_1_instruction_master_translator:uav_write -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_1_instruction_master_translator:uav_read -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_1_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_1_instruction_master_translator:uav_readdata
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_1_instruction_master_translator:uav_debugaccess -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_1_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_1_instruction_master_translator:uav_byteenable -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_1_instruction_master_translator:uav_readdatavalid
	wire         cpu_1_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_1_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_1_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_1_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_1_data_master_translator:uav_burstcount -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_1_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_1_data_master_translator:uav_writedata -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_1_data_master_translator_avalon_universal_master_0_address;                                     // cpu_1_data_master_translator:uav_address -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_1_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_1_data_master_translator:uav_lock -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_1_data_master_translator_avalon_universal_master_0_write;                                       // cpu_1_data_master_translator:uav_write -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_1_data_master_translator_avalon_universal_master_0_read;                                        // cpu_1_data_master_translator:uav_read -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_1_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_1_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_1_data_master_translator:uav_readdata
	wire         cpu_1_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_1_data_master_translator:uav_debugaccess -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_1_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_1_data_master_translator:uav_byteenable -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_1_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_1_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_1_data_master_translator:uav_readdatavalid
	wire         cpu_0_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_0_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_0_data_master_translator:uav_burstcount -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_0_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_0_data_master_translator:uav_writedata -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [13:0] cpu_0_data_master_translator_avalon_universal_master_0_address;                                     // cpu_0_data_master_translator:uav_address -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_0_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_0_data_master_translator:uav_lock -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_0_data_master_translator_avalon_universal_master_0_write;                                       // cpu_0_data_master_translator:uav_write -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_0_data_master_translator_avalon_universal_master_0_read;                                        // cpu_0_data_master_translator:uav_read -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_0_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_data_master_translator:uav_readdata
	wire         cpu_0_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_0_data_master_translator:uav_debugaccess -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_0_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_0_data_master_translator:uav_byteenable -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_data_master_translator:uav_readdatavalid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_0_jtag_debug_module_translator:uav_waitrequest -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_0_jtag_debug_module_translator:uav_writedata
	wire  [13:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_0_jtag_debug_module_translator:uav_address
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_0_jtag_debug_module_translator:uav_write
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_0_jtag_debug_module_translator:uav_lock
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_0_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_0_jtag_debug_module_translator:uav_readdata -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_0_jtag_debug_module_translator:uav_readdatavalid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_0_jtag_debug_module_translator:uav_byteenable
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // ins_mem_0_s1_translator:uav_waitrequest -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ins_mem_0_s1_translator:uav_burstcount
	wire  [31:0] ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ins_mem_0_s1_translator:uav_writedata
	wire  [13:0] ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> ins_mem_0_s1_translator:uav_address
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> ins_mem_0_s1_translator:uav_write
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ins_mem_0_s1_translator:uav_lock
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> ins_mem_0_s1_translator:uav_read
	wire  [31:0] ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // ins_mem_0_s1_translator:uav_readdata -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // ins_mem_0_s1_translator:uav_readdatavalid -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ins_mem_0_s1_translator:uav_debugaccess
	wire   [3:0] ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ins_mem_0_s1_translator:uav_byteenable
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // atob_0_in_translator:uav_waitrequest -> atob_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atob_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // atob_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> atob_0_in_translator:uav_burstcount
	wire  [31:0] atob_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // atob_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> atob_0_in_translator:uav_writedata
	wire  [13:0] atob_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // atob_0_in_translator_avalon_universal_slave_0_agent:m0_address -> atob_0_in_translator:uav_address
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // atob_0_in_translator_avalon_universal_slave_0_agent:m0_write -> atob_0_in_translator:uav_write
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // atob_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> atob_0_in_translator:uav_lock
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // atob_0_in_translator_avalon_universal_slave_0_agent:m0_read -> atob_0_in_translator:uav_read
	wire  [31:0] atob_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // atob_0_in_translator:uav_readdata -> atob_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // atob_0_in_translator:uav_readdatavalid -> atob_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // atob_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atob_0_in_translator:uav_debugaccess
	wire   [3:0] atob_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // atob_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> atob_0_in_translator:uav_byteenable
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // atob_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // atob_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // atob_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // atob_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atob_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atob_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atob_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atob_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atob_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // atob_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // atob_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atob_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atob_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // atob_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atob_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // atob_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atob_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // atob_0_in_csr_translator:uav_waitrequest -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> atob_0_in_csr_translator:uav_burstcount
	wire  [31:0] atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> atob_0_in_csr_translator:uav_writedata
	wire  [13:0] atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> atob_0_in_csr_translator:uav_address
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> atob_0_in_csr_translator:uav_write
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> atob_0_in_csr_translator:uav_lock
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> atob_0_in_csr_translator:uav_read
	wire  [31:0] atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // atob_0_in_csr_translator:uav_readdata -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // atob_0_in_csr_translator:uav_readdatavalid -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atob_0_in_csr_translator:uav_debugaccess
	wire   [3:0] atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // atob_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> atob_0_in_csr_translator:uav_byteenable
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atob_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // atob_0_out_translator:uav_waitrequest -> atob_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atob_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // atob_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> atob_0_out_translator:uav_burstcount
	wire  [31:0] atob_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // atob_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> atob_0_out_translator:uav_writedata
	wire  [13:0] atob_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // atob_0_out_translator_avalon_universal_slave_0_agent:m0_address -> atob_0_out_translator:uav_address
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // atob_0_out_translator_avalon_universal_slave_0_agent:m0_write -> atob_0_out_translator:uav_write
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // atob_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> atob_0_out_translator:uav_lock
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // atob_0_out_translator_avalon_universal_slave_0_agent:m0_read -> atob_0_out_translator:uav_read
	wire  [31:0] atob_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // atob_0_out_translator:uav_readdata -> atob_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // atob_0_out_translator:uav_readdatavalid -> atob_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // atob_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atob_0_out_translator:uav_debugaccess
	wire   [3:0] atob_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // atob_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> atob_0_out_translator:uav_byteenable
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // atob_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // atob_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // atob_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // atob_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atob_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atob_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atob_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atob_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atob_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // atob_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // atob_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atob_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atob_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // atob_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atob_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // atob_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atob_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // atob_1_in_translator:uav_waitrequest -> atob_1_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atob_1_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // atob_1_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> atob_1_in_translator:uav_burstcount
	wire  [31:0] atob_1_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // atob_1_in_translator_avalon_universal_slave_0_agent:m0_writedata -> atob_1_in_translator:uav_writedata
	wire  [13:0] atob_1_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // atob_1_in_translator_avalon_universal_slave_0_agent:m0_address -> atob_1_in_translator:uav_address
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // atob_1_in_translator_avalon_universal_slave_0_agent:m0_write -> atob_1_in_translator:uav_write
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // atob_1_in_translator_avalon_universal_slave_0_agent:m0_lock -> atob_1_in_translator:uav_lock
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // atob_1_in_translator_avalon_universal_slave_0_agent:m0_read -> atob_1_in_translator:uav_read
	wire  [31:0] atob_1_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // atob_1_in_translator:uav_readdata -> atob_1_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // atob_1_in_translator:uav_readdatavalid -> atob_1_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // atob_1_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atob_1_in_translator:uav_debugaccess
	wire   [3:0] atob_1_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // atob_1_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> atob_1_in_translator:uav_byteenable
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // atob_1_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // atob_1_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // atob_1_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // atob_1_in_translator_avalon_universal_slave_0_agent:rf_source_data -> atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atob_1_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atob_1_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atob_1_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atob_1_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atob_1_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // atob_1_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // atob_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atob_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atob_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // atob_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atob_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // atob_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atob_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // atob_1_in_csr_translator:uav_waitrequest -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> atob_1_in_csr_translator:uav_burstcount
	wire  [31:0] atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> atob_1_in_csr_translator:uav_writedata
	wire  [13:0] atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> atob_1_in_csr_translator:uav_address
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> atob_1_in_csr_translator:uav_write
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> atob_1_in_csr_translator:uav_lock
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> atob_1_in_csr_translator:uav_read
	wire  [31:0] atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // atob_1_in_csr_translator:uav_readdata -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // atob_1_in_csr_translator:uav_readdatavalid -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atob_1_in_csr_translator:uav_debugaccess
	wire   [3:0] atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // atob_1_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> atob_1_in_csr_translator:uav_byteenable
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atob_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // atob_1_out_translator:uav_waitrequest -> atob_1_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atob_1_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // atob_1_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> atob_1_out_translator:uav_burstcount
	wire  [31:0] atob_1_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // atob_1_out_translator_avalon_universal_slave_0_agent:m0_writedata -> atob_1_out_translator:uav_writedata
	wire  [13:0] atob_1_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // atob_1_out_translator_avalon_universal_slave_0_agent:m0_address -> atob_1_out_translator:uav_address
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // atob_1_out_translator_avalon_universal_slave_0_agent:m0_write -> atob_1_out_translator:uav_write
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // atob_1_out_translator_avalon_universal_slave_0_agent:m0_lock -> atob_1_out_translator:uav_lock
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // atob_1_out_translator_avalon_universal_slave_0_agent:m0_read -> atob_1_out_translator:uav_read
	wire  [31:0] atob_1_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // atob_1_out_translator:uav_readdata -> atob_1_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // atob_1_out_translator:uav_readdatavalid -> atob_1_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // atob_1_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atob_1_out_translator:uav_debugaccess
	wire   [3:0] atob_1_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // atob_1_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> atob_1_out_translator:uav_byteenable
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // atob_1_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // atob_1_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // atob_1_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // atob_1_out_translator_avalon_universal_slave_0_agent:rf_source_data -> atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atob_1_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atob_1_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atob_1_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atob_1_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atob_1_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // atob_1_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // atob_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atob_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atob_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // atob_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atob_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // atob_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atob_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // atob_2_in_translator:uav_waitrequest -> atob_2_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atob_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // atob_2_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> atob_2_in_translator:uav_burstcount
	wire  [31:0] atob_2_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // atob_2_in_translator_avalon_universal_slave_0_agent:m0_writedata -> atob_2_in_translator:uav_writedata
	wire  [13:0] atob_2_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // atob_2_in_translator_avalon_universal_slave_0_agent:m0_address -> atob_2_in_translator:uav_address
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // atob_2_in_translator_avalon_universal_slave_0_agent:m0_write -> atob_2_in_translator:uav_write
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // atob_2_in_translator_avalon_universal_slave_0_agent:m0_lock -> atob_2_in_translator:uav_lock
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // atob_2_in_translator_avalon_universal_slave_0_agent:m0_read -> atob_2_in_translator:uav_read
	wire  [31:0] atob_2_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // atob_2_in_translator:uav_readdata -> atob_2_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // atob_2_in_translator:uav_readdatavalid -> atob_2_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // atob_2_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atob_2_in_translator:uav_debugaccess
	wire   [3:0] atob_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // atob_2_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> atob_2_in_translator:uav_byteenable
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // atob_2_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // atob_2_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // atob_2_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // atob_2_in_translator_avalon_universal_slave_0_agent:rf_source_data -> atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atob_2_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atob_2_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atob_2_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atob_2_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atob_2_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // atob_2_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // atob_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atob_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atob_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // atob_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atob_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // atob_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atob_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // atob_2_in_csr_translator:uav_waitrequest -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> atob_2_in_csr_translator:uav_burstcount
	wire  [31:0] atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> atob_2_in_csr_translator:uav_writedata
	wire  [13:0] atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> atob_2_in_csr_translator:uav_address
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> atob_2_in_csr_translator:uav_write
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> atob_2_in_csr_translator:uav_lock
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> atob_2_in_csr_translator:uav_read
	wire  [31:0] atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // atob_2_in_csr_translator:uav_readdata -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // atob_2_in_csr_translator:uav_readdatavalid -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atob_2_in_csr_translator:uav_debugaccess
	wire   [3:0] atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // atob_2_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> atob_2_in_csr_translator:uav_byteenable
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atob_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // atob_2_out_translator:uav_waitrequest -> atob_2_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atob_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // atob_2_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> atob_2_out_translator:uav_burstcount
	wire  [31:0] atob_2_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // atob_2_out_translator_avalon_universal_slave_0_agent:m0_writedata -> atob_2_out_translator:uav_writedata
	wire  [13:0] atob_2_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // atob_2_out_translator_avalon_universal_slave_0_agent:m0_address -> atob_2_out_translator:uav_address
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // atob_2_out_translator_avalon_universal_slave_0_agent:m0_write -> atob_2_out_translator:uav_write
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // atob_2_out_translator_avalon_universal_slave_0_agent:m0_lock -> atob_2_out_translator:uav_lock
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // atob_2_out_translator_avalon_universal_slave_0_agent:m0_read -> atob_2_out_translator:uav_read
	wire  [31:0] atob_2_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // atob_2_out_translator:uav_readdata -> atob_2_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // atob_2_out_translator:uav_readdatavalid -> atob_2_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // atob_2_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atob_2_out_translator:uav_debugaccess
	wire   [3:0] atob_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // atob_2_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> atob_2_out_translator:uav_byteenable
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // atob_2_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // atob_2_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // atob_2_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // atob_2_out_translator_avalon_universal_slave_0_agent:rf_source_data -> atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atob_2_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atob_2_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atob_2_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atob_2_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atob_2_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // atob_2_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // atob_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atob_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atob_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // atob_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atob_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // atob_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atob_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // atod_0_in_translator:uav_waitrequest -> atod_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atod_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // atod_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> atod_0_in_translator:uav_burstcount
	wire  [31:0] atod_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // atod_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> atod_0_in_translator:uav_writedata
	wire  [13:0] atod_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // atod_0_in_translator_avalon_universal_slave_0_agent:m0_address -> atod_0_in_translator:uav_address
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // atod_0_in_translator_avalon_universal_slave_0_agent:m0_write -> atod_0_in_translator:uav_write
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // atod_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> atod_0_in_translator:uav_lock
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // atod_0_in_translator_avalon_universal_slave_0_agent:m0_read -> atod_0_in_translator:uav_read
	wire  [31:0] atod_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // atod_0_in_translator:uav_readdata -> atod_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // atod_0_in_translator:uav_readdatavalid -> atod_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // atod_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atod_0_in_translator:uav_debugaccess
	wire   [3:0] atod_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // atod_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> atod_0_in_translator:uav_byteenable
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // atod_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // atod_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // atod_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // atod_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atod_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // atod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // atod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // atod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // atod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // atod_0_out_translator:uav_waitrequest -> atod_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atod_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // atod_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> atod_0_out_translator:uav_burstcount
	wire  [31:0] atod_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // atod_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> atod_0_out_translator:uav_writedata
	wire  [13:0] atod_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // atod_0_out_translator_avalon_universal_slave_0_agent:m0_address -> atod_0_out_translator:uav_address
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // atod_0_out_translator_avalon_universal_slave_0_agent:m0_write -> atod_0_out_translator:uav_write
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // atod_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> atod_0_out_translator:uav_lock
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // atod_0_out_translator_avalon_universal_slave_0_agent:m0_read -> atod_0_out_translator:uav_read
	wire  [31:0] atod_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // atod_0_out_translator:uav_readdata -> atod_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // atod_0_out_translator:uav_readdatavalid -> atod_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // atod_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atod_0_out_translator:uav_debugaccess
	wire   [3:0] atod_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // atod_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> atod_0_out_translator:uav_byteenable
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // atod_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // atod_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // atod_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // atod_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atod_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // atod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // atod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // atod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // atod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // atod_0_in_csr_translator:uav_waitrequest -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> atod_0_in_csr_translator:uav_burstcount
	wire  [31:0] atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> atod_0_in_csr_translator:uav_writedata
	wire  [13:0] atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> atod_0_in_csr_translator:uav_address
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> atod_0_in_csr_translator:uav_write
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> atod_0_in_csr_translator:uav_lock
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> atod_0_in_csr_translator:uav_read
	wire  [31:0] atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // atod_0_in_csr_translator:uav_readdata -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // atod_0_in_csr_translator:uav_readdatavalid -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atod_0_in_csr_translator:uav_debugaccess
	wire   [3:0] atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // atod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> atod_0_in_csr_translator:uav_byteenable
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // atoe_0_in_translator:uav_waitrequest -> atoe_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atoe_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // atoe_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> atoe_0_in_translator:uav_burstcount
	wire  [31:0] atoe_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // atoe_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> atoe_0_in_translator:uav_writedata
	wire  [13:0] atoe_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // atoe_0_in_translator_avalon_universal_slave_0_agent:m0_address -> atoe_0_in_translator:uav_address
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // atoe_0_in_translator_avalon_universal_slave_0_agent:m0_write -> atoe_0_in_translator:uav_write
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // atoe_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> atoe_0_in_translator:uav_lock
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // atoe_0_in_translator_avalon_universal_slave_0_agent:m0_read -> atoe_0_in_translator:uav_read
	wire  [31:0] atoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // atoe_0_in_translator:uav_readdata -> atoe_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // atoe_0_in_translator:uav_readdatavalid -> atoe_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // atoe_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atoe_0_in_translator:uav_debugaccess
	wire   [3:0] atoe_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // atoe_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> atoe_0_in_translator:uav_byteenable
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // atoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // atoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // atoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // atoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // atoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // atoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // atoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // atoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // atoe_0_out_translator:uav_waitrequest -> atoe_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atoe_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // atoe_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> atoe_0_out_translator:uav_burstcount
	wire  [31:0] atoe_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // atoe_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> atoe_0_out_translator:uav_writedata
	wire  [13:0] atoe_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // atoe_0_out_translator_avalon_universal_slave_0_agent:m0_address -> atoe_0_out_translator:uav_address
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // atoe_0_out_translator_avalon_universal_slave_0_agent:m0_write -> atoe_0_out_translator:uav_write
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // atoe_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> atoe_0_out_translator:uav_lock
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // atoe_0_out_translator_avalon_universal_slave_0_agent:m0_read -> atoe_0_out_translator:uav_read
	wire  [31:0] atoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // atoe_0_out_translator:uav_readdata -> atoe_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // atoe_0_out_translator:uav_readdatavalid -> atoe_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // atoe_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atoe_0_out_translator:uav_debugaccess
	wire   [3:0] atoe_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // atoe_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> atoe_0_out_translator:uav_byteenable
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // atoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // atoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // atoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // atoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // atoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // atoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // atoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // atoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // atoe_0_in_csr_translator:uav_waitrequest -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> atoe_0_in_csr_translator:uav_burstcount
	wire  [31:0] atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> atoe_0_in_csr_translator:uav_writedata
	wire  [13:0] atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> atoe_0_in_csr_translator:uav_address
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> atoe_0_in_csr_translator:uav_write
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> atoe_0_in_csr_translator:uav_lock
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> atoe_0_in_csr_translator:uav_read
	wire  [31:0] atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // atoe_0_in_csr_translator:uav_readdata -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // atoe_0_in_csr_translator:uav_readdatavalid -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atoe_0_in_csr_translator:uav_debugaccess
	wire   [3:0] atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> atoe_0_in_csr_translator:uav_byteenable
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // atof_0_in_translator:uav_waitrequest -> atof_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atof_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // atof_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> atof_0_in_translator:uav_burstcount
	wire  [31:0] atof_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // atof_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> atof_0_in_translator:uav_writedata
	wire  [13:0] atof_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // atof_0_in_translator_avalon_universal_slave_0_agent:m0_address -> atof_0_in_translator:uav_address
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // atof_0_in_translator_avalon_universal_slave_0_agent:m0_write -> atof_0_in_translator:uav_write
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // atof_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> atof_0_in_translator:uav_lock
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // atof_0_in_translator_avalon_universal_slave_0_agent:m0_read -> atof_0_in_translator:uav_read
	wire  [31:0] atof_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // atof_0_in_translator:uav_readdata -> atof_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // atof_0_in_translator:uav_readdatavalid -> atof_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // atof_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atof_0_in_translator:uav_debugaccess
	wire   [3:0] atof_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // atof_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> atof_0_in_translator:uav_byteenable
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // atof_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // atof_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // atof_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // atof_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atof_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // atof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // atof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // atof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // atof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // atof_0_in_csr_translator:uav_waitrequest -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> atof_0_in_csr_translator:uav_burstcount
	wire  [31:0] atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> atof_0_in_csr_translator:uav_writedata
	wire  [13:0] atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> atof_0_in_csr_translator:uav_address
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> atof_0_in_csr_translator:uav_write
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> atof_0_in_csr_translator:uav_lock
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> atof_0_in_csr_translator:uav_read
	wire  [31:0] atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // atof_0_in_csr_translator:uav_readdata -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // atof_0_in_csr_translator:uav_readdatavalid -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atof_0_in_csr_translator:uav_debugaccess
	wire   [3:0] atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // atof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> atof_0_in_csr_translator:uav_byteenable
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // atof_0_out_translator:uav_waitrequest -> atof_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] atof_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // atof_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> atof_0_out_translator:uav_burstcount
	wire  [31:0] atof_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // atof_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> atof_0_out_translator:uav_writedata
	wire  [13:0] atof_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // atof_0_out_translator_avalon_universal_slave_0_agent:m0_address -> atof_0_out_translator:uav_address
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // atof_0_out_translator_avalon_universal_slave_0_agent:m0_write -> atof_0_out_translator:uav_write
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // atof_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> atof_0_out_translator:uav_lock
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // atof_0_out_translator_avalon_universal_slave_0_agent:m0_read -> atof_0_out_translator:uav_read
	wire  [31:0] atof_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // atof_0_out_translator:uav_readdata -> atof_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // atof_0_out_translator:uav_readdatavalid -> atof_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // atof_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> atof_0_out_translator:uav_debugaccess
	wire   [3:0] atof_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // atof_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> atof_0_out_translator:uav_byteenable
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // atof_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // atof_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // atof_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // atof_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> atof_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> atof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> atof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> atof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> atof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // atof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // atof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> atof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] atof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // atof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> atof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // atof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> atof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // ins_mem_5_s1_translator:uav_waitrequest -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ins_mem_5_s1_translator:uav_burstcount
	wire  [31:0] ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ins_mem_5_s1_translator:uav_writedata
	wire  [13:0] ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_address -> ins_mem_5_s1_translator:uav_address
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_write -> ins_mem_5_s1_translator:uav_write
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ins_mem_5_s1_translator:uav_lock
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_read -> ins_mem_5_s1_translator:uav_read
	wire  [31:0] ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // ins_mem_5_s1_translator:uav_readdata -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // ins_mem_5_s1_translator:uav_readdatavalid -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ins_mem_5_s1_translator:uav_debugaccess
	wire   [3:0] ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ins_mem_5_s1_translator:uav_byteenable
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_5_jtag_debug_module_translator:uav_waitrequest -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_5_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_5_jtag_debug_module_translator:uav_writedata
	wire  [13:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_5_jtag_debug_module_translator:uav_address
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_5_jtag_debug_module_translator:uav_write
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_5_jtag_debug_module_translator:uav_lock
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_5_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_5_jtag_debug_module_translator:uav_readdata -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_5_jtag_debug_module_translator:uav_readdatavalid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_5_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_5_jtag_debug_module_translator:uav_byteenable
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // etof_0_in_translator:uav_waitrequest -> etof_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] etof_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // etof_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> etof_0_in_translator:uav_burstcount
	wire  [31:0] etof_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // etof_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> etof_0_in_translator:uav_writedata
	wire  [13:0] etof_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // etof_0_in_translator_avalon_universal_slave_0_agent:m0_address -> etof_0_in_translator:uav_address
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // etof_0_in_translator_avalon_universal_slave_0_agent:m0_write -> etof_0_in_translator:uav_write
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // etof_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> etof_0_in_translator:uav_lock
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // etof_0_in_translator_avalon_universal_slave_0_agent:m0_read -> etof_0_in_translator:uav_read
	wire  [31:0] etof_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // etof_0_in_translator:uav_readdata -> etof_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // etof_0_in_translator:uav_readdatavalid -> etof_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // etof_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> etof_0_in_translator:uav_debugaccess
	wire   [3:0] etof_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // etof_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> etof_0_in_translator:uav_byteenable
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // etof_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // etof_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // etof_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // etof_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> etof_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> etof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> etof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> etof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> etof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // etof_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // etof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> etof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] etof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // etof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> etof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // etof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> etof_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // etof_0_in_csr_translator:uav_waitrequest -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> etof_0_in_csr_translator:uav_burstcount
	wire  [31:0] etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> etof_0_in_csr_translator:uav_writedata
	wire  [13:0] etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> etof_0_in_csr_translator:uav_address
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> etof_0_in_csr_translator:uav_write
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> etof_0_in_csr_translator:uav_lock
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> etof_0_in_csr_translator:uav_read
	wire  [31:0] etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // etof_0_in_csr_translator:uav_readdata -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // etof_0_in_csr_translator:uav_readdatavalid -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> etof_0_in_csr_translator:uav_debugaccess
	wire   [3:0] etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // etof_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> etof_0_in_csr_translator:uav_byteenable
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] etof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // etof_0_out_translator:uav_waitrequest -> etof_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] etof_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // etof_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> etof_0_out_translator:uav_burstcount
	wire  [31:0] etof_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // etof_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> etof_0_out_translator:uav_writedata
	wire  [13:0] etof_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // etof_0_out_translator_avalon_universal_slave_0_agent:m0_address -> etof_0_out_translator:uav_address
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // etof_0_out_translator_avalon_universal_slave_0_agent:m0_write -> etof_0_out_translator:uav_write
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // etof_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> etof_0_out_translator:uav_lock
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // etof_0_out_translator_avalon_universal_slave_0_agent:m0_read -> etof_0_out_translator:uav_read
	wire  [31:0] etof_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // etof_0_out_translator:uav_readdata -> etof_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // etof_0_out_translator:uav_readdatavalid -> etof_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // etof_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> etof_0_out_translator:uav_debugaccess
	wire   [3:0] etof_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // etof_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> etof_0_out_translator:uav_byteenable
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // etof_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // etof_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // etof_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // etof_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> etof_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> etof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> etof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> etof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> etof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // etof_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // etof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> etof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] etof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // etof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> etof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // etof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> etof_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // data_mem_5_s1_translator:uav_waitrequest -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> data_mem_5_s1_translator:uav_burstcount
	wire  [31:0] data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> data_mem_5_s1_translator:uav_writedata
	wire  [13:0] data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_address -> data_mem_5_s1_translator:uav_address
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_write -> data_mem_5_s1_translator:uav_write
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> data_mem_5_s1_translator:uav_lock
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_read -> data_mem_5_s1_translator:uav_read
	wire  [31:0] data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // data_mem_5_s1_translator:uav_readdata -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // data_mem_5_s1_translator:uav_readdatavalid -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> data_mem_5_s1_translator:uav_debugaccess
	wire   [3:0] data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // data_mem_5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> data_mem_5_s1_translator:uav_byteenable
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_5_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_5_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_5_avalon_jtag_slave_translator:uav_writedata
	wire  [13:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_5_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_5_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_5_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_5_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_5_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_5_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_5_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_5_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_5_s1_translator:uav_waitrequest -> timer_5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_5_s1_translator:uav_burstcount
	wire  [31:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_5_s1_translator:uav_writedata
	wire  [13:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_5_s1_translator:uav_address
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_5_s1_translator:uav_write
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_5_s1_translator:uav_lock
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_5_s1_translator:uav_read
	wire  [31:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_5_s1_translator:uav_readdata -> timer_5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_5_s1_translator:uav_readdatavalid -> timer_5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_5_s1_translator:uav_debugaccess
	wire   [3:0] timer_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_5_s1_translator:uav_byteenable
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // high_scale_timer_5_s1_translator:uav_waitrequest -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_scale_timer_5_s1_translator:uav_burstcount
	wire  [31:0] high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_scale_timer_5_s1_translator:uav_writedata
	wire  [13:0] high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_scale_timer_5_s1_translator:uav_address
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_scale_timer_5_s1_translator:uav_write
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_scale_timer_5_s1_translator:uav_lock
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_scale_timer_5_s1_translator:uav_read
	wire  [31:0] high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // high_scale_timer_5_s1_translator:uav_readdata -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // high_scale_timer_5_s1_translator:uav_readdatavalid -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_scale_timer_5_s1_translator:uav_debugaccess
	wire   [3:0] high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_scale_timer_5_s1_translator:uav_byteenable
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // ins_mem_4_s1_translator:uav_waitrequest -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ins_mem_4_s1_translator:uav_burstcount
	wire  [31:0] ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ins_mem_4_s1_translator:uav_writedata
	wire  [13:0] ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> ins_mem_4_s1_translator:uav_address
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> ins_mem_4_s1_translator:uav_write
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ins_mem_4_s1_translator:uav_lock
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> ins_mem_4_s1_translator:uav_read
	wire  [31:0] ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // ins_mem_4_s1_translator:uav_readdata -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // ins_mem_4_s1_translator:uav_readdatavalid -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ins_mem_4_s1_translator:uav_debugaccess
	wire   [3:0] ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ins_mem_4_s1_translator:uav_byteenable
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_4_jtag_debug_module_translator:uav_waitrequest -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_4_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_4_jtag_debug_module_translator:uav_writedata
	wire  [13:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_4_jtag_debug_module_translator:uav_address
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_4_jtag_debug_module_translator:uav_write
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_4_jtag_debug_module_translator:uav_lock
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_4_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_4_jtag_debug_module_translator:uav_readdata -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_4_jtag_debug_module_translator:uav_readdatavalid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_4_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_4_jtag_debug_module_translator:uav_byteenable
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // dtoe_0_in_translator:uav_waitrequest -> dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> dtoe_0_in_translator:uav_burstcount
	wire  [31:0] dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> dtoe_0_in_translator:uav_writedata
	wire  [13:0] dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_address -> dtoe_0_in_translator:uav_address
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_write -> dtoe_0_in_translator:uav_write
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> dtoe_0_in_translator:uav_lock
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_read -> dtoe_0_in_translator:uav_read
	wire  [31:0] dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // dtoe_0_in_translator:uav_readdata -> dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // dtoe_0_in_translator:uav_readdatavalid -> dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dtoe_0_in_translator:uav_debugaccess
	wire   [3:0] dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // dtoe_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> dtoe_0_in_translator:uav_byteenable
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // dtoe_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // dtoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dtoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] dtoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // dtoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dtoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // dtoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dtoe_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // dtoe_0_in_csr_translator:uav_waitrequest -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> dtoe_0_in_csr_translator:uav_burstcount
	wire  [31:0] dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> dtoe_0_in_csr_translator:uav_writedata
	wire  [13:0] dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> dtoe_0_in_csr_translator:uav_address
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> dtoe_0_in_csr_translator:uav_write
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> dtoe_0_in_csr_translator:uav_lock
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> dtoe_0_in_csr_translator:uav_read
	wire  [31:0] dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // dtoe_0_in_csr_translator:uav_readdata -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // dtoe_0_in_csr_translator:uav_readdatavalid -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dtoe_0_in_csr_translator:uav_debugaccess
	wire   [3:0] dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> dtoe_0_in_csr_translator:uav_byteenable
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // dtoe_0_out_translator:uav_waitrequest -> dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> dtoe_0_out_translator:uav_burstcount
	wire  [31:0] dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> dtoe_0_out_translator:uav_writedata
	wire  [13:0] dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_address -> dtoe_0_out_translator:uav_address
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_write -> dtoe_0_out_translator:uav_write
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> dtoe_0_out_translator:uav_lock
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_read -> dtoe_0_out_translator:uav_read
	wire  [31:0] dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // dtoe_0_out_translator:uav_readdata -> dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // dtoe_0_out_translator:uav_readdatavalid -> dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dtoe_0_out_translator:uav_debugaccess
	wire   [3:0] dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // dtoe_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> dtoe_0_out_translator:uav_byteenable
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // dtoe_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // dtoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dtoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] dtoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // dtoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dtoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // dtoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dtoe_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // data_mem_4_s1_translator:uav_waitrequest -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> data_mem_4_s1_translator:uav_burstcount
	wire  [31:0] data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> data_mem_4_s1_translator:uav_writedata
	wire  [13:0] data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> data_mem_4_s1_translator:uav_address
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> data_mem_4_s1_translator:uav_write
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> data_mem_4_s1_translator:uav_lock
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> data_mem_4_s1_translator:uav_read
	wire  [31:0] data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // data_mem_4_s1_translator:uav_readdata -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // data_mem_4_s1_translator:uav_readdatavalid -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> data_mem_4_s1_translator:uav_debugaccess
	wire   [3:0] data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // data_mem_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> data_mem_4_s1_translator:uav_byteenable
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_4_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_4_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_4_avalon_jtag_slave_translator:uav_writedata
	wire  [13:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_4_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_4_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_4_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_4_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_4_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_4_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_4_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_4_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_4_s1_translator:uav_waitrequest -> timer_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_4_s1_translator:uav_burstcount
	wire  [31:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_4_s1_translator:uav_writedata
	wire  [13:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_4_s1_translator:uav_address
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_4_s1_translator:uav_write
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_4_s1_translator:uav_lock
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_4_s1_translator:uav_read
	wire  [31:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_4_s1_translator:uav_readdata -> timer_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_4_s1_translator:uav_readdatavalid -> timer_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_4_s1_translator:uav_debugaccess
	wire   [3:0] timer_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_4_s1_translator:uav_byteenable
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // high_scale_timer_4_s1_translator:uav_waitrequest -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_scale_timer_4_s1_translator:uav_burstcount
	wire  [31:0] high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_scale_timer_4_s1_translator:uav_writedata
	wire  [13:0] high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_scale_timer_4_s1_translator:uav_address
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_scale_timer_4_s1_translator:uav_write
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_scale_timer_4_s1_translator:uav_lock
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_scale_timer_4_s1_translator:uav_read
	wire  [31:0] high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // high_scale_timer_4_s1_translator:uav_readdata -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // high_scale_timer_4_s1_translator:uav_readdatavalid -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_scale_timer_4_s1_translator:uav_debugaccess
	wire   [3:0] high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_scale_timer_4_s1_translator:uav_byteenable
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // ins_mem_3_s1_translator:uav_waitrequest -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ins_mem_3_s1_translator:uav_burstcount
	wire  [31:0] ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ins_mem_3_s1_translator:uav_writedata
	wire  [13:0] ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> ins_mem_3_s1_translator:uav_address
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> ins_mem_3_s1_translator:uav_write
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ins_mem_3_s1_translator:uav_lock
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> ins_mem_3_s1_translator:uav_read
	wire  [31:0] ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // ins_mem_3_s1_translator:uav_readdata -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // ins_mem_3_s1_translator:uav_readdatavalid -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ins_mem_3_s1_translator:uav_debugaccess
	wire   [3:0] ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ins_mem_3_s1_translator:uav_byteenable
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_3_jtag_debug_module_translator:uav_waitrequest -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_3_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_3_jtag_debug_module_translator:uav_writedata
	wire  [13:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_3_jtag_debug_module_translator:uav_address
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_3_jtag_debug_module_translator:uav_write
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_3_jtag_debug_module_translator:uav_lock
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_3_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_3_jtag_debug_module_translator:uav_readdata -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_3_jtag_debug_module_translator:uav_readdatavalid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_3_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_3_jtag_debug_module_translator:uav_byteenable
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // ctod_0_in_translator:uav_waitrequest -> ctod_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ctod_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // ctod_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> ctod_0_in_translator:uav_burstcount
	wire  [31:0] ctod_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // ctod_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> ctod_0_in_translator:uav_writedata
	wire  [13:0] ctod_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // ctod_0_in_translator_avalon_universal_slave_0_agent:m0_address -> ctod_0_in_translator:uav_address
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // ctod_0_in_translator_avalon_universal_slave_0_agent:m0_write -> ctod_0_in_translator:uav_write
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // ctod_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> ctod_0_in_translator:uav_lock
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // ctod_0_in_translator_avalon_universal_slave_0_agent:m0_read -> ctod_0_in_translator:uav_read
	wire  [31:0] ctod_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // ctod_0_in_translator:uav_readdata -> ctod_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // ctod_0_in_translator:uav_readdatavalid -> ctod_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // ctod_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ctod_0_in_translator:uav_debugaccess
	wire   [3:0] ctod_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // ctod_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> ctod_0_in_translator:uav_byteenable
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // ctod_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // ctod_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // ctod_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // ctod_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ctod_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ctod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ctod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ctod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ctod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // ctod_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // ctod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ctod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ctod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // ctod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ctod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // ctod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ctod_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // ctod_0_in_csr_translator:uav_waitrequest -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> ctod_0_in_csr_translator:uav_burstcount
	wire  [31:0] ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> ctod_0_in_csr_translator:uav_writedata
	wire  [13:0] ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> ctod_0_in_csr_translator:uav_address
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> ctod_0_in_csr_translator:uav_write
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> ctod_0_in_csr_translator:uav_lock
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> ctod_0_in_csr_translator:uav_read
	wire  [31:0] ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // ctod_0_in_csr_translator:uav_readdata -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // ctod_0_in_csr_translator:uav_readdatavalid -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ctod_0_in_csr_translator:uav_debugaccess
	wire   [3:0] ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> ctod_0_in_csr_translator:uav_byteenable
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // ctod_0_out_translator:uav_waitrequest -> ctod_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ctod_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // ctod_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> ctod_0_out_translator:uav_burstcount
	wire  [31:0] ctod_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // ctod_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> ctod_0_out_translator:uav_writedata
	wire  [13:0] ctod_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // ctod_0_out_translator_avalon_universal_slave_0_agent:m0_address -> ctod_0_out_translator:uav_address
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // ctod_0_out_translator_avalon_universal_slave_0_agent:m0_write -> ctod_0_out_translator:uav_write
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // ctod_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> ctod_0_out_translator:uav_lock
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // ctod_0_out_translator_avalon_universal_slave_0_agent:m0_read -> ctod_0_out_translator:uav_read
	wire  [31:0] ctod_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // ctod_0_out_translator:uav_readdata -> ctod_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // ctod_0_out_translator:uav_readdatavalid -> ctod_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // ctod_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ctod_0_out_translator:uav_debugaccess
	wire   [3:0] ctod_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // ctod_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> ctod_0_out_translator:uav_byteenable
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // ctod_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // ctod_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // ctod_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // ctod_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ctod_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ctod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ctod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ctod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ctod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // ctod_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // ctod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ctod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ctod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // ctod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ctod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // ctod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ctod_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // data_mem_3_s1_translator:uav_waitrequest -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> data_mem_3_s1_translator:uav_burstcount
	wire  [31:0] data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> data_mem_3_s1_translator:uav_writedata
	wire  [13:0] data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> data_mem_3_s1_translator:uav_address
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> data_mem_3_s1_translator:uav_write
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> data_mem_3_s1_translator:uav_lock
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> data_mem_3_s1_translator:uav_read
	wire  [31:0] data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // data_mem_3_s1_translator:uav_readdata -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // data_mem_3_s1_translator:uav_readdatavalid -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> data_mem_3_s1_translator:uav_debugaccess
	wire   [3:0] data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // data_mem_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> data_mem_3_s1_translator:uav_byteenable
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_3_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_3_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_3_avalon_jtag_slave_translator:uav_writedata
	wire  [13:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_3_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_3_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_3_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_3_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_3_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_3_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_3_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_3_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_3_s1_translator:uav_waitrequest -> timer_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_3_s1_translator:uav_burstcount
	wire  [31:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_3_s1_translator:uav_writedata
	wire  [13:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_3_s1_translator:uav_address
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_3_s1_translator:uav_write
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_3_s1_translator:uav_lock
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_3_s1_translator:uav_read
	wire  [31:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_3_s1_translator:uav_readdata -> timer_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_3_s1_translator:uav_readdatavalid -> timer_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_3_s1_translator:uav_debugaccess
	wire   [3:0] timer_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_3_s1_translator:uav_byteenable
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // high_scale_timer_3_s1_translator:uav_waitrequest -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_scale_timer_3_s1_translator:uav_burstcount
	wire  [31:0] high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_scale_timer_3_s1_translator:uav_writedata
	wire  [13:0] high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_scale_timer_3_s1_translator:uav_address
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_scale_timer_3_s1_translator:uav_write
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_scale_timer_3_s1_translator:uav_lock
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_scale_timer_3_s1_translator:uav_read
	wire  [31:0] high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // high_scale_timer_3_s1_translator:uav_readdata -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // high_scale_timer_3_s1_translator:uav_readdatavalid -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_scale_timer_3_s1_translator:uav_debugaccess
	wire   [3:0] high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_scale_timer_3_s1_translator:uav_byteenable
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // data_mem_2_s1_translator:uav_waitrequest -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> data_mem_2_s1_translator:uav_burstcount
	wire  [31:0] data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> data_mem_2_s1_translator:uav_writedata
	wire  [13:0] data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> data_mem_2_s1_translator:uav_address
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> data_mem_2_s1_translator:uav_write
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> data_mem_2_s1_translator:uav_lock
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> data_mem_2_s1_translator:uav_read
	wire  [31:0] data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // data_mem_2_s1_translator:uav_readdata -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // data_mem_2_s1_translator:uav_readdatavalid -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> data_mem_2_s1_translator:uav_debugaccess
	wire   [3:0] data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // data_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> data_mem_2_s1_translator:uav_byteenable
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_2_jtag_debug_module_translator:uav_waitrequest -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_2_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_2_jtag_debug_module_translator:uav_writedata
	wire  [13:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_2_jtag_debug_module_translator:uav_address
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_2_jtag_debug_module_translator:uav_write
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_2_jtag_debug_module_translator:uav_lock
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_2_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_2_jtag_debug_module_translator:uav_readdata -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_2_jtag_debug_module_translator:uav_readdatavalid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_2_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_2_jtag_debug_module_translator:uav_byteenable
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_2_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_2_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_2_avalon_jtag_slave_translator:uav_writedata
	wire  [13:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_2_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_2_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_2_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_2_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_2_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_2_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_2_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_2_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_2_s1_translator:uav_waitrequest -> timer_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_2_s1_translator:uav_burstcount
	wire  [31:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_2_s1_translator:uav_writedata
	wire  [13:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_2_s1_translator:uav_address
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_2_s1_translator:uav_write
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_2_s1_translator:uav_lock
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_2_s1_translator:uav_read
	wire  [31:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_2_s1_translator:uav_readdata -> timer_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_2_s1_translator:uav_readdatavalid -> timer_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_2_s1_translator:uav_debugaccess
	wire   [3:0] timer_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_2_s1_translator:uav_byteenable
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // high_scale_timer_2_s1_translator:uav_waitrequest -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_scale_timer_2_s1_translator:uav_burstcount
	wire  [31:0] high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_scale_timer_2_s1_translator:uav_writedata
	wire  [13:0] high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_scale_timer_2_s1_translator:uav_address
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_scale_timer_2_s1_translator:uav_write
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_scale_timer_2_s1_translator:uav_lock
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_scale_timer_2_s1_translator:uav_read
	wire  [31:0] high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // high_scale_timer_2_s1_translator:uav_readdata -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // high_scale_timer_2_s1_translator:uav_readdatavalid -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_scale_timer_2_s1_translator:uav_debugaccess
	wire   [3:0] high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_scale_timer_2_s1_translator:uav_byteenable
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // btoc_0_in_translator:uav_waitrequest -> btoc_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] btoc_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // btoc_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> btoc_0_in_translator:uav_burstcount
	wire  [31:0] btoc_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // btoc_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> btoc_0_in_translator:uav_writedata
	wire  [13:0] btoc_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                     // btoc_0_in_translator_avalon_universal_slave_0_agent:m0_address -> btoc_0_in_translator:uav_address
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                       // btoc_0_in_translator_avalon_universal_slave_0_agent:m0_write -> btoc_0_in_translator:uav_write
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                        // btoc_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> btoc_0_in_translator:uav_lock
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                        // btoc_0_in_translator_avalon_universal_slave_0_agent:m0_read -> btoc_0_in_translator:uav_read
	wire  [31:0] btoc_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // btoc_0_in_translator:uav_readdata -> btoc_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // btoc_0_in_translator:uav_readdatavalid -> btoc_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // btoc_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> btoc_0_in_translator:uav_debugaccess
	wire   [3:0] btoc_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // btoc_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> btoc_0_in_translator:uav_byteenable
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // btoc_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // btoc_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // btoc_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // btoc_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> btoc_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> btoc_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> btoc_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> btoc_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> btoc_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // btoc_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // btoc_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> btoc_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] btoc_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // btoc_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> btoc_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // btoc_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> btoc_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // btoc_0_out_translator:uav_waitrequest -> btoc_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] btoc_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // btoc_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> btoc_0_out_translator:uav_burstcount
	wire  [31:0] btoc_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // btoc_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> btoc_0_out_translator:uav_writedata
	wire  [13:0] btoc_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                    // btoc_0_out_translator_avalon_universal_slave_0_agent:m0_address -> btoc_0_out_translator:uav_address
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                      // btoc_0_out_translator_avalon_universal_slave_0_agent:m0_write -> btoc_0_out_translator:uav_write
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                       // btoc_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> btoc_0_out_translator:uav_lock
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                       // btoc_0_out_translator_avalon_universal_slave_0_agent:m0_read -> btoc_0_out_translator:uav_read
	wire  [31:0] btoc_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // btoc_0_out_translator:uav_readdata -> btoc_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // btoc_0_out_translator:uav_readdatavalid -> btoc_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // btoc_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> btoc_0_out_translator:uav_debugaccess
	wire   [3:0] btoc_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // btoc_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> btoc_0_out_translator:uav_byteenable
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // btoc_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // btoc_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // btoc_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                // btoc_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> btoc_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> btoc_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> btoc_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> btoc_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> btoc_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // btoc_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // btoc_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> btoc_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] btoc_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // btoc_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> btoc_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // btoc_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> btoc_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // btoc_0_in_csr_translator:uav_waitrequest -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> btoc_0_in_csr_translator:uav_burstcount
	wire  [31:0] btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> btoc_0_in_csr_translator:uav_writedata
	wire  [13:0] btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> btoc_0_in_csr_translator:uav_address
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> btoc_0_in_csr_translator:uav_write
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> btoc_0_in_csr_translator:uav_lock
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> btoc_0_in_csr_translator:uav_read
	wire  [31:0] btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // btoc_0_in_csr_translator:uav_readdata -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // btoc_0_in_csr_translator:uav_readdatavalid -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> btoc_0_in_csr_translator:uav_debugaccess
	wire   [3:0] btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> btoc_0_in_csr_translator:uav_byteenable
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // ins_mem_2_s1_translator:uav_waitrequest -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ins_mem_2_s1_translator:uav_burstcount
	wire  [31:0] ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ins_mem_2_s1_translator:uav_writedata
	wire  [13:0] ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> ins_mem_2_s1_translator:uav_address
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> ins_mem_2_s1_translator:uav_write
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ins_mem_2_s1_translator:uav_lock
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> ins_mem_2_s1_translator:uav_read
	wire  [31:0] ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // ins_mem_2_s1_translator:uav_readdata -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // ins_mem_2_s1_translator:uav_readdatavalid -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ins_mem_2_s1_translator:uav_debugaccess
	wire   [3:0] ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ins_mem_2_s1_translator:uav_byteenable
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // ins_mem_1_s1_translator:uav_waitrequest -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ins_mem_1_s1_translator:uav_burstcount
	wire  [31:0] ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ins_mem_1_s1_translator:uav_writedata
	wire  [13:0] ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> ins_mem_1_s1_translator:uav_address
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> ins_mem_1_s1_translator:uav_write
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ins_mem_1_s1_translator:uav_lock
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> ins_mem_1_s1_translator:uav_read
	wire  [31:0] ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // ins_mem_1_s1_translator:uav_readdata -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // ins_mem_1_s1_translator:uav_readdatavalid -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ins_mem_1_s1_translator:uav_debugaccess
	wire   [3:0] ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ins_mem_1_s1_translator:uav_byteenable
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_1_jtag_debug_module_translator:uav_waitrequest -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_1_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_1_jtag_debug_module_translator:uav_writedata
	wire  [13:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_1_jtag_debug_module_translator:uav_address
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_1_jtag_debug_module_translator:uav_write
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_1_jtag_debug_module_translator:uav_lock
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_1_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_1_jtag_debug_module_translator:uav_readdata -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_1_jtag_debug_module_translator:uav_readdatavalid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_1_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_1_jtag_debug_module_translator:uav_byteenable
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // data_mem_1_s1_translator:uav_waitrequest -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> data_mem_1_s1_translator:uav_burstcount
	wire  [31:0] data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> data_mem_1_s1_translator:uav_writedata
	wire  [13:0] data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> data_mem_1_s1_translator:uav_address
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> data_mem_1_s1_translator:uav_write
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> data_mem_1_s1_translator:uav_lock
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> data_mem_1_s1_translator:uav_read
	wire  [31:0] data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // data_mem_1_s1_translator:uav_readdata -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // data_mem_1_s1_translator:uav_readdatavalid -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> data_mem_1_s1_translator:uav_debugaccess
	wire   [3:0] data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // data_mem_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> data_mem_1_s1_translator:uav_byteenable
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_1_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_1_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_1_avalon_jtag_slave_translator:uav_writedata
	wire  [13:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_1_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_1_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_1_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_1_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_1_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_1_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_1_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_1_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	wire  [13:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	wire   [3:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // high_scale_timer_1_s1_translator:uav_waitrequest -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_scale_timer_1_s1_translator:uav_burstcount
	wire  [31:0] high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_scale_timer_1_s1_translator:uav_writedata
	wire  [13:0] high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_scale_timer_1_s1_translator:uav_address
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_scale_timer_1_s1_translator:uav_write
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_scale_timer_1_s1_translator:uav_lock
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_scale_timer_1_s1_translator:uav_read
	wire  [31:0] high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // high_scale_timer_1_s1_translator:uav_readdata -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // high_scale_timer_1_s1_translator:uav_readdatavalid -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_scale_timer_1_s1_translator:uav_debugaccess
	wire   [3:0] high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_scale_timer_1_s1_translator:uav_byteenable
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // data_mem_0_s1_translator:uav_waitrequest -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> data_mem_0_s1_translator:uav_burstcount
	wire  [31:0] data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> data_mem_0_s1_translator:uav_writedata
	wire  [13:0] data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> data_mem_0_s1_translator:uav_address
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> data_mem_0_s1_translator:uav_write
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> data_mem_0_s1_translator:uav_lock
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> data_mem_0_s1_translator:uav_read
	wire  [31:0] data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // data_mem_0_s1_translator:uav_readdata -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // data_mem_0_s1_translator:uav_readdatavalid -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> data_mem_0_s1_translator:uav_debugaccess
	wire   [3:0] data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // data_mem_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> data_mem_0_s1_translator:uav_byteenable
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [13:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [13:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // high_scale_timer_0_s1_translator:uav_waitrequest -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_scale_timer_0_s1_translator:uav_burstcount
	wire  [31:0] high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_scale_timer_0_s1_translator:uav_writedata
	wire  [13:0] high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_scale_timer_0_s1_translator:uav_address
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_scale_timer_0_s1_translator:uav_write
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_scale_timer_0_s1_translator:uav_lock
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_scale_timer_0_s1_translator:uav_read
	wire  [31:0] high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // high_scale_timer_0_s1_translator:uav_readdata -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // high_scale_timer_0_s1_translator:uav_readdatavalid -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_scale_timer_0_s1_translator:uav_debugaccess
	wire   [3:0] high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_scale_timer_0_s1_translator:uav_byteenable
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [94:0] cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router:sink_ready -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [94:0] cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_001:sink_ready -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire         cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire         cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [94:0] cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire         cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_002:sink_ready -> cpu_5_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [94:0] cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire         cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_003:sink_ready -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire         cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire         cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [94:0] cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire         cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_004:sink_ready -> cpu_4_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [94:0] cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire         cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_005:sink_ready -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire         cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire         cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire  [94:0] cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire         cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_006:sink_ready -> cpu_3_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	wire         cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	wire         cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	wire  [94:0] cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	wire         cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_007:sink_ready -> cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_008:sink_endofpacket
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_008:sink_valid
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_008:sink_startofpacket
	wire  [94:0] cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_008:sink_data
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_008:sink_ready -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_009:sink_endofpacket
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_009:sink_valid
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_009:sink_startofpacket
	wire  [94:0] cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_009:sink_data
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_009:sink_ready -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_010:sink_endofpacket
	wire         cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_010:sink_valid
	wire         cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_010:sink_startofpacket
	wire  [94:0] cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_010:sink_data
	wire         cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_010:sink_ready -> cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_011:sink_endofpacket
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_011:sink_valid
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_011:sink_startofpacket
	wire  [94:0] cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_011:sink_data
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_011:sink_ready -> cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [94:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router:sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [94:0] ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_001:sink_ready -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // atob_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // atob_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // atob_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [94:0] atob_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // atob_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         atob_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_002:sink_ready -> atob_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [94:0] atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // atob_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_003:sink_ready -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // atob_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // atob_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // atob_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [94:0] atob_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // atob_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         atob_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_004:sink_ready -> atob_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // atob_1_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // atob_1_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // atob_1_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [94:0] atob_1_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // atob_1_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         atob_1_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_005:sink_ready -> atob_1_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [94:0] atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // atob_1_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_006:sink_ready -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // atob_1_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // atob_1_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // atob_1_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [94:0] atob_1_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // atob_1_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         atob_1_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_007:sink_ready -> atob_1_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // atob_2_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // atob_2_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // atob_2_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [94:0] atob_2_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // atob_2_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         atob_2_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_008:sink_ready -> atob_2_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [94:0] atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // atob_2_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_009:sink_ready -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // atob_2_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // atob_2_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // atob_2_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [94:0] atob_2_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // atob_2_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         atob_2_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_010:sink_ready -> atob_2_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // atod_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // atod_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // atod_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [94:0] atod_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // atod_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         atod_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_011:sink_ready -> atod_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // atod_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // atod_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // atod_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [94:0] atod_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // atod_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         atod_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_012:sink_ready -> atod_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [94:0] atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // atod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_013:sink_ready -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // atoe_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // atoe_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // atoe_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [94:0] atoe_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // atoe_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire         atoe_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_014:sink_ready -> atoe_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // atoe_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // atoe_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // atoe_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [94:0] atoe_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // atoe_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire         atoe_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_015:sink_ready -> atoe_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [94:0] atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire         atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_016:sink_ready -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // atof_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // atof_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // atof_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [94:0] atof_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // atof_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire         atof_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_017:sink_ready -> atof_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [94:0] atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // atof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire         atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_018:sink_ready -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // atof_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // atof_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // atof_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [94:0] atof_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // atof_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire         atof_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_019:sink_ready -> atof_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [94:0] ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire         ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_020:sink_ready -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [94:0] cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire         cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_021:sink_ready -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // etof_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // etof_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // etof_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [94:0] etof_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // etof_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire         etof_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_022:sink_ready -> etof_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire  [94:0] etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // etof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire         etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_023:sink_ready -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // etof_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // etof_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // etof_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire  [94:0] etof_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // etof_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire         etof_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_024:sink_ready -> etof_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire  [94:0] data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // data_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire         data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_025:sink_ready -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire  [94:0] jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire         jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_026:sink_ready -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire  [94:0] timer_5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire         timer_5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_027:sink_ready -> timer_5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire  [94:0] high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire         high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_028:sink_ready -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire  [94:0] ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire         ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_029:sink_ready -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire  [94:0] cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire         cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_030:sink_ready -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // dtoe_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // dtoe_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // dtoe_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	wire  [94:0] dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // dtoe_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	wire         dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_031:sink_ready -> dtoe_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	wire  [94:0] dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	wire         dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_032:sink_ready -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // dtoe_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_033:sink_endofpacket
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // dtoe_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_033:sink_valid
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // dtoe_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_033:sink_startofpacket
	wire  [94:0] dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // dtoe_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_033:sink_data
	wire         dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_033:sink_ready -> dtoe_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_034:sink_endofpacket
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_034:sink_valid
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_034:sink_startofpacket
	wire  [94:0] data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // data_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_034:sink_data
	wire         data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_034:sink_ready -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_035:sink_endofpacket
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_035:sink_valid
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_035:sink_startofpacket
	wire  [94:0] jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_035:sink_data
	wire         jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_035:sink_ready -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_036:sink_endofpacket
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_036:sink_valid
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_036:sink_startofpacket
	wire  [94:0] timer_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_036:sink_data
	wire         timer_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_036:sink_ready -> timer_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_037:sink_endofpacket
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_037:sink_valid
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_037:sink_startofpacket
	wire  [94:0] high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_037:sink_data
	wire         high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_037:sink_ready -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_038:sink_endofpacket
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_038:sink_valid
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_038:sink_startofpacket
	wire  [94:0] ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_038:sink_data
	wire         ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_038:sink_ready -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_039:sink_endofpacket
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_039:sink_valid
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_039:sink_startofpacket
	wire  [94:0] cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_039:sink_data
	wire         cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_039:sink_ready -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // ctod_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_040:sink_endofpacket
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // ctod_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_040:sink_valid
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // ctod_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_040:sink_startofpacket
	wire  [94:0] ctod_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // ctod_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_040:sink_data
	wire         ctod_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_040:sink_ready -> ctod_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_041:sink_endofpacket
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_041:sink_valid
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_041:sink_startofpacket
	wire  [94:0] ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_041:sink_data
	wire         ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_041:sink_ready -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // ctod_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_042:sink_endofpacket
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // ctod_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_042:sink_valid
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // ctod_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_042:sink_startofpacket
	wire  [94:0] ctod_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // ctod_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_042:sink_data
	wire         ctod_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_042:sink_ready -> ctod_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_043:sink_endofpacket
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_043:sink_valid
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_043:sink_startofpacket
	wire  [94:0] data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // data_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_043:sink_data
	wire         data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_043:sink_ready -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_044:sink_endofpacket
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_044:sink_valid
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_044:sink_startofpacket
	wire  [94:0] jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_044:sink_data
	wire         jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_044:sink_ready -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_045:sink_endofpacket
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_045:sink_valid
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_045:sink_startofpacket
	wire  [94:0] timer_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_045:sink_data
	wire         timer_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_045:sink_ready -> timer_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_046:sink_endofpacket
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_046:sink_valid
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_046:sink_startofpacket
	wire  [94:0] high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_046:sink_data
	wire         high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_046:sink_ready -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_047:sink_endofpacket
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_047:sink_valid
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_047:sink_startofpacket
	wire  [94:0] data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // data_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_047:sink_data
	wire         data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_047:sink_ready -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_048:sink_endofpacket
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_048:sink_valid
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_048:sink_startofpacket
	wire  [94:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_048:sink_data
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_048:sink_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_049:sink_endofpacket
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_049:sink_valid
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_049:sink_startofpacket
	wire  [94:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_049:sink_data
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_049:sink_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_050:sink_endofpacket
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_050:sink_valid
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_050:sink_startofpacket
	wire  [94:0] timer_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_050:sink_data
	wire         timer_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_050:sink_ready -> timer_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_051:sink_endofpacket
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_051:sink_valid
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_051:sink_startofpacket
	wire  [94:0] high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_051:sink_data
	wire         high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_051:sink_ready -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // btoc_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_052:sink_endofpacket
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                       // btoc_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_052:sink_valid
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // btoc_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_052:sink_startofpacket
	wire  [94:0] btoc_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                        // btoc_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_052:sink_data
	wire         btoc_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_052:sink_ready -> btoc_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // btoc_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_053:sink_endofpacket
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                      // btoc_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_053:sink_valid
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // btoc_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_053:sink_startofpacket
	wire  [94:0] btoc_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                       // btoc_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_053:sink_data
	wire         btoc_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_053:sink_ready -> btoc_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_054:sink_endofpacket
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_054:sink_valid
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_054:sink_startofpacket
	wire  [94:0] btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_054:sink_data
	wire         btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_054:sink_ready -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_055:sink_endofpacket
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_055:sink_valid
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_055:sink_startofpacket
	wire  [94:0] ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_055:sink_data
	wire         ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_055:sink_ready -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_056:sink_endofpacket
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_056:sink_valid
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_056:sink_startofpacket
	wire  [94:0] ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_056:sink_data
	wire         ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_056:sink_ready -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_057:sink_endofpacket
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_057:sink_valid
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_057:sink_startofpacket
	wire  [94:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_057:sink_data
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_057:sink_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_058:sink_endofpacket
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_058:sink_valid
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_058:sink_startofpacket
	wire  [94:0] data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // data_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_058:sink_data
	wire         data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_058:sink_ready -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_059:sink_endofpacket
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_059:sink_valid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_059:sink_startofpacket
	wire  [94:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_059:sink_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_059:sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_060:sink_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_060:sink_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_060:sink_startofpacket
	wire  [94:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_060:sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_060:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_061:sink_endofpacket
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_061:sink_valid
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_061:sink_startofpacket
	wire  [94:0] high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_061:sink_data
	wire         high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_061:sink_ready -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_062:sink_endofpacket
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_062:sink_valid
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_062:sink_startofpacket
	wire  [94:0] data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // data_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_062:sink_data
	wire         data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_062:sink_ready -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_063:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_063:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_063:sink_startofpacket
	wire  [94:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_063:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_063:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_064:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_064:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_064:sink_startofpacket
	wire  [94:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_064:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_064:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_065:sink_endofpacket
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_065:sink_valid
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_065:sink_startofpacket
	wire  [94:0] high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_065:sink_data
	wire         high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_065:sink_ready -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                        // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                              // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                      // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [94:0] addr_router_src_data;                                                                               // addr_router:src_data -> limiter:cmd_sink_data
	wire  [65:0] addr_router_src_channel;                                                                            // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                              // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                        // limiter:rsp_src_endofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                              // limiter:rsp_src_valid -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                      // limiter:rsp_src_startofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] limiter_rsp_src_data;                                                                               // limiter:rsp_src_data -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] limiter_rsp_src_channel;                                                                            // limiter:rsp_src_channel -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                              // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                    // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                          // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                  // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [94:0] addr_router_001_src_data;                                                                           // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire  [65:0] addr_router_001_src_channel;                                                                        // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                          // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                    // limiter_001:rsp_src_endofpacket -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                          // limiter_001:rsp_src_valid -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                  // limiter_001:rsp_src_startofpacket -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] limiter_001_rsp_src_data;                                                                           // limiter_001:rsp_src_data -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] limiter_001_rsp_src_channel;                                                                        // limiter_001:rsp_src_channel -> cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                          // cpu_5_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         addr_router_003_src_endofpacket;                                                                    // addr_router_003:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire         addr_router_003_src_valid;                                                                          // addr_router_003:src_valid -> limiter_002:cmd_sink_valid
	wire         addr_router_003_src_startofpacket;                                                                  // addr_router_003:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire  [94:0] addr_router_003_src_data;                                                                           // addr_router_003:src_data -> limiter_002:cmd_sink_data
	wire  [65:0] addr_router_003_src_channel;                                                                        // addr_router_003:src_channel -> limiter_002:cmd_sink_channel
	wire         addr_router_003_src_ready;                                                                          // limiter_002:cmd_sink_ready -> addr_router_003:src_ready
	wire         limiter_002_rsp_src_endofpacket;                                                                    // limiter_002:rsp_src_endofpacket -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_002_rsp_src_valid;                                                                          // limiter_002:rsp_src_valid -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_002_rsp_src_startofpacket;                                                                  // limiter_002:rsp_src_startofpacket -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] limiter_002_rsp_src_data;                                                                           // limiter_002:rsp_src_data -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] limiter_002_rsp_src_channel;                                                                        // limiter_002:rsp_src_channel -> cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_002_rsp_src_ready;                                                                          // cpu_4_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire         addr_router_005_src_endofpacket;                                                                    // addr_router_005:src_endofpacket -> limiter_003:cmd_sink_endofpacket
	wire         addr_router_005_src_valid;                                                                          // addr_router_005:src_valid -> limiter_003:cmd_sink_valid
	wire         addr_router_005_src_startofpacket;                                                                  // addr_router_005:src_startofpacket -> limiter_003:cmd_sink_startofpacket
	wire  [94:0] addr_router_005_src_data;                                                                           // addr_router_005:src_data -> limiter_003:cmd_sink_data
	wire  [65:0] addr_router_005_src_channel;                                                                        // addr_router_005:src_channel -> limiter_003:cmd_sink_channel
	wire         addr_router_005_src_ready;                                                                          // limiter_003:cmd_sink_ready -> addr_router_005:src_ready
	wire         limiter_003_rsp_src_endofpacket;                                                                    // limiter_003:rsp_src_endofpacket -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_003_rsp_src_valid;                                                                          // limiter_003:rsp_src_valid -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_003_rsp_src_startofpacket;                                                                  // limiter_003:rsp_src_startofpacket -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] limiter_003_rsp_src_data;                                                                           // limiter_003:rsp_src_data -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] limiter_003_rsp_src_channel;                                                                        // limiter_003:rsp_src_channel -> cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_003_rsp_src_ready;                                                                          // cpu_3_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_003:rsp_src_ready
	wire         addr_router_008_src_endofpacket;                                                                    // addr_router_008:src_endofpacket -> limiter_004:cmd_sink_endofpacket
	wire         addr_router_008_src_valid;                                                                          // addr_router_008:src_valid -> limiter_004:cmd_sink_valid
	wire         addr_router_008_src_startofpacket;                                                                  // addr_router_008:src_startofpacket -> limiter_004:cmd_sink_startofpacket
	wire  [94:0] addr_router_008_src_data;                                                                           // addr_router_008:src_data -> limiter_004:cmd_sink_data
	wire  [65:0] addr_router_008_src_channel;                                                                        // addr_router_008:src_channel -> limiter_004:cmd_sink_channel
	wire         addr_router_008_src_ready;                                                                          // limiter_004:cmd_sink_ready -> addr_router_008:src_ready
	wire         limiter_004_rsp_src_endofpacket;                                                                    // limiter_004:rsp_src_endofpacket -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_004_rsp_src_valid;                                                                          // limiter_004:rsp_src_valid -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_004_rsp_src_startofpacket;                                                                  // limiter_004:rsp_src_startofpacket -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] limiter_004_rsp_src_data;                                                                           // limiter_004:rsp_src_data -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] limiter_004_rsp_src_channel;                                                                        // limiter_004:rsp_src_channel -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_004_rsp_src_ready;                                                                          // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_004:rsp_src_ready
	wire         addr_router_009_src_endofpacket;                                                                    // addr_router_009:src_endofpacket -> limiter_005:cmd_sink_endofpacket
	wire         addr_router_009_src_valid;                                                                          // addr_router_009:src_valid -> limiter_005:cmd_sink_valid
	wire         addr_router_009_src_startofpacket;                                                                  // addr_router_009:src_startofpacket -> limiter_005:cmd_sink_startofpacket
	wire  [94:0] addr_router_009_src_data;                                                                           // addr_router_009:src_data -> limiter_005:cmd_sink_data
	wire  [65:0] addr_router_009_src_channel;                                                                        // addr_router_009:src_channel -> limiter_005:cmd_sink_channel
	wire         addr_router_009_src_ready;                                                                          // limiter_005:cmd_sink_ready -> addr_router_009:src_ready
	wire         limiter_005_rsp_src_endofpacket;                                                                    // limiter_005:rsp_src_endofpacket -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_005_rsp_src_valid;                                                                          // limiter_005:rsp_src_valid -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_005_rsp_src_startofpacket;                                                                  // limiter_005:rsp_src_startofpacket -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] limiter_005_rsp_src_data;                                                                           // limiter_005:rsp_src_data -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] limiter_005_rsp_src_channel;                                                                        // limiter_005:rsp_src_channel -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_005_rsp_src_ready;                                                                          // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_005:rsp_src_ready
	wire         rst_controller_reset_out_reset;                                                                     // rst_controller:reset_out -> [addr_router:reset, addr_router_011:reset, cmd_xbar_demux:reset, cmd_xbar_demux_011:reset, cmd_xbar_mux:reset, cpu_0:reset_n, cpu_0_data_master_translator:reset, cpu_0_data_master_translator_avalon_universal_master_0_agent:reset, cpu_0_instruction_master_translator:reset, cpu_0_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_0_jtag_debug_module_translator:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, data_mem_0:reset, data_mem_0_s1_translator:reset, data_mem_0_s1_translator_avalon_universal_slave_0_agent:reset, data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, high_scale_timer_0:reset_n, high_scale_timer_0_s1_translator:reset, high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:reset, high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_062:reset, id_router_063:reset, id_router_064:reset, id_router_065:reset, ins_mem_0:reset, ins_mem_0_s1_translator:reset, ins_mem_0_s1_translator_avalon_universal_slave_0_agent:reset, ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_062:reset, rsp_xbar_demux_063:reset, rsp_xbar_demux_064:reset, rsp_xbar_demux_065:reset, rsp_xbar_mux:reset, rsp_xbar_mux_011:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cpu_0_jtag_debug_module_reset_reset;                                                                // cpu_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_007:reset_in1, rst_controller_012:reset_in2, rst_controller_013:reset_in1, rst_controller_014:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                                                 // rst_controller_001:reset_out -> [data_mem_1:reset, data_mem_1_s1_translator:reset, data_mem_1_s1_translator_avalon_universal_slave_0_agent:reset, data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, high_scale_timer_1:reset_n, high_scale_timer_1_s1_translator:reset, high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:reset, high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_056:reset, id_router_058:reset, id_router_059:reset, id_router_060:reset, id_router_061:reset, ins_mem_1:reset, ins_mem_1_s1_translator:reset, ins_mem_1_s1_translator_avalon_universal_slave_0_agent:reset, ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, jtag_uart_1:rst_n, jtag_uart_1_avalon_jtag_slave_translator:reset, jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_056:reset, rsp_xbar_demux_058:reset, rsp_xbar_demux_059:reset, rsp_xbar_demux_060:reset, rsp_xbar_demux_061:reset, timer_1:reset_n, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cpu_1_jtag_debug_module_reset_reset;                                                                // cpu_1:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in1, rst_controller_007:reset_in2, rst_controller_008:reset_in2]
	wire         rst_controller_002_reset_out_reset;                                                                 // rst_controller_002:reset_out -> [addr_router_009:reset, addr_router_010:reset, cmd_xbar_demux_009:reset, cmd_xbar_demux_010:reset, cmd_xbar_mux_057:reset, cpu_1:reset_n, cpu_1_data_master_translator:reset, cpu_1_data_master_translator_avalon_universal_master_0_agent:reset, cpu_1_instruction_master_translator:reset, cpu_1_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_1_jtag_debug_module_translator:reset, cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_057:reset, irq_mapper_001:reset, limiter_005:reset, rsp_xbar_demux_057:reset, rsp_xbar_mux_009:reset, rsp_xbar_mux_010:reset]
	wire         rst_controller_003_reset_out_reset;                                                                 // rst_controller_003:reset_out -> [addr_router_007:reset, addr_router_008:reset, cmd_xbar_demux_007:reset, cmd_xbar_demux_008:reset, cmd_xbar_mux_048:reset, cpu_2:reset_n, cpu_2_data_master_translator:reset, cpu_2_data_master_translator_avalon_universal_master_0_agent:reset, cpu_2_instruction_master_translator:reset, cpu_2_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_2_jtag_debug_module_translator:reset, cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, data_mem_2:reset, data_mem_2_s1_translator:reset, data_mem_2_s1_translator_avalon_universal_slave_0_agent:reset, data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, high_scale_timer_2:reset_n, high_scale_timer_2_s1_translator:reset, high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:reset, high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_047:reset, id_router_048:reset, id_router_049:reset, id_router_050:reset, id_router_051:reset, id_router_055:reset, ins_mem_2:reset, ins_mem_2_s1_translator:reset, ins_mem_2_s1_translator_avalon_universal_slave_0_agent:reset, ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, irq_mapper_002:reset, jtag_uart_2:rst_n, jtag_uart_2_avalon_jtag_slave_translator:reset, jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_004:reset, rsp_xbar_demux_047:reset, rsp_xbar_demux_048:reset, rsp_xbar_demux_049:reset, rsp_xbar_demux_050:reset, rsp_xbar_demux_051:reset, rsp_xbar_demux_055:reset, rsp_xbar_mux_007:reset, rsp_xbar_mux_008:reset, timer_2:reset_n, timer_2_s1_translator:reset, timer_2_s1_translator_avalon_universal_slave_0_agent:reset, timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cpu_2_jtag_debug_module_reset_reset;                                                                // cpu_2:jtag_debug_module_resetrequest -> [rst_controller_003:reset_in1, rst_controller_008:reset_in1, rst_controller_009:reset_in2]
	wire         rst_controller_004_reset_out_reset;                                                                 // rst_controller_004:reset_out -> [addr_router_005:reset, addr_router_006:reset, cmd_xbar_demux_005:reset, cmd_xbar_demux_006:reset, cmd_xbar_mux_039:reset, cpu_3:reset_n, cpu_3_data_master_translator:reset, cpu_3_data_master_translator_avalon_universal_master_0_agent:reset, cpu_3_instruction_master_translator:reset, cpu_3_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_3_jtag_debug_module_translator:reset, cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, data_mem_3:reset, data_mem_3_s1_translator:reset, data_mem_3_s1_translator_avalon_universal_slave_0_agent:reset, data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, high_scale_timer_3:reset_n, high_scale_timer_3_s1_translator:reset, high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:reset, high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_038:reset, id_router_039:reset, id_router_043:reset, id_router_044:reset, id_router_045:reset, id_router_046:reset, ins_mem_3:reset, ins_mem_3_s1_translator:reset, ins_mem_3_s1_translator_avalon_universal_slave_0_agent:reset, ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, irq_mapper_003:reset, jtag_uart_3:rst_n, jtag_uart_3_avalon_jtag_slave_translator:reset, jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_003:reset, rsp_xbar_demux_038:reset, rsp_xbar_demux_039:reset, rsp_xbar_demux_043:reset, rsp_xbar_demux_044:reset, rsp_xbar_demux_045:reset, rsp_xbar_demux_046:reset, rsp_xbar_mux_005:reset, rsp_xbar_mux_006:reset, timer_3:reset_n, timer_3_s1_translator:reset, timer_3_s1_translator_avalon_universal_slave_0_agent:reset, timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cpu_3_jtag_debug_module_reset_reset;                                                                // cpu_3:jtag_debug_module_resetrequest -> [rst_controller_004:reset_in1, rst_controller_009:reset_in1, rst_controller_010:reset_in1, rst_controller_013:reset_in2]
	wire         rst_controller_005_reset_out_reset;                                                                 // rst_controller_005:reset_out -> [addr_router_003:reset, addr_router_004:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux_030:reset, cpu_4:reset_n, cpu_4_data_master_translator:reset, cpu_4_data_master_translator_avalon_universal_master_0_agent:reset, cpu_4_instruction_master_translator:reset, cpu_4_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_4_jtag_debug_module_translator:reset, cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, data_mem_4:reset, data_mem_4_s1_translator:reset, data_mem_4_s1_translator_avalon_universal_slave_0_agent:reset, data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, high_scale_timer_4:reset_n, high_scale_timer_4_s1_translator:reset, high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:reset, high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_029:reset, id_router_030:reset, id_router_034:reset, id_router_035:reset, id_router_036:reset, id_router_037:reset, ins_mem_4:reset, ins_mem_4_s1_translator:reset, ins_mem_4_s1_translator_avalon_universal_slave_0_agent:reset, ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, irq_mapper_004:reset, jtag_uart_4:rst_n, jtag_uart_4_avalon_jtag_slave_translator:reset, jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_002:reset, rsp_xbar_demux_029:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_034:reset, rsp_xbar_demux_035:reset, rsp_xbar_demux_036:reset, rsp_xbar_demux_037:reset, rsp_xbar_mux_003:reset, rsp_xbar_mux_004:reset, timer_4:reset_n, timer_4_s1_translator:reset, timer_4_s1_translator_avalon_universal_slave_0_agent:reset, timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cpu_4_jtag_debug_module_reset_reset;                                                                // cpu_4:jtag_debug_module_resetrequest -> [rst_controller_005:reset_in1, rst_controller_010:reset_in2, rst_controller_011:reset_in1, rst_controller_014:reset_in2]
	wire         rst_controller_006_reset_out_reset;                                                                 // rst_controller_006:reset_out -> [addr_router_001:reset, addr_router_002:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_mux_021:reset, cpu_5:reset_n, cpu_5_data_master_translator:reset, cpu_5_data_master_translator_avalon_universal_master_0_agent:reset, cpu_5_instruction_master_translator:reset, cpu_5_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_5_jtag_debug_module_translator:reset, cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, data_mem_5:reset, data_mem_5_s1_translator:reset, data_mem_5_s1_translator_avalon_universal_slave_0_agent:reset, data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, high_scale_timer_5:reset_n, high_scale_timer_5_s1_translator:reset, high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:reset, high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_020:reset, id_router_021:reset, id_router_025:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, ins_mem_5:reset, ins_mem_5_s1_translator:reset, ins_mem_5_s1_translator_avalon_universal_slave_0_agent:reset, ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, irq_mapper_005:reset, jtag_uart_5:rst_n, jtag_uart_5_avalon_jtag_slave_translator:reset, jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_001:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, timer_5:reset_n, timer_5_s1_translator:reset, timer_5_s1_translator_avalon_universal_slave_0_agent:reset, timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cpu_5_jtag_debug_module_reset_reset;                                                                // cpu_5:jtag_debug_module_resetrequest -> [rst_controller_006:reset_in1, rst_controller_011:reset_in2, rst_controller_012:reset_in1]
	wire         rst_controller_007_reset_out_reset;                                                                 // rst_controller_007:reset_out -> [atob_0:reset_n, atob_0_in_csr_translator:reset, atob_0_in_csr_translator_avalon_universal_slave_0_agent:reset, atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atob_0_in_translator:reset, atob_0_in_translator_avalon_universal_slave_0_agent:reset, atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atob_0_out_translator:reset, atob_0_out_translator_avalon_universal_slave_0_agent:reset, atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atob_1:reset_n, atob_1_in_csr_translator:reset, atob_1_in_csr_translator_avalon_universal_slave_0_agent:reset, atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atob_1_in_translator:reset, atob_1_in_translator_avalon_universal_slave_0_agent:reset, atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atob_1_out_translator:reset, atob_1_out_translator_avalon_universal_slave_0_agent:reset, atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atob_2:reset_n, atob_2_in_csr_translator:reset, atob_2_in_csr_translator_avalon_universal_slave_0_agent:reset, atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atob_2_in_translator:reset, atob_2_in_translator_avalon_universal_slave_0_agent:reset, atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atob_2_out_translator:reset, atob_2_out_translator_avalon_universal_slave_0_agent:reset, atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, cmd_xbar_mux_010:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset]
	wire         rst_controller_008_reset_out_reset;                                                                 // rst_controller_008:reset_out -> [btoc_0:reset_n, btoc_0_in_csr_translator:reset, btoc_0_in_csr_translator_avalon_universal_slave_0_agent:reset, btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, btoc_0_in_translator:reset, btoc_0_in_translator_avalon_universal_slave_0_agent:reset, btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, btoc_0_out_translator:reset, btoc_0_out_translator_avalon_universal_slave_0_agent:reset, btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_052:reset, cmd_xbar_mux_053:reset, cmd_xbar_mux_054:reset, id_router_052:reset, id_router_053:reset, id_router_054:reset, rsp_xbar_demux_052:reset, rsp_xbar_demux_053:reset, rsp_xbar_demux_054:reset]
	wire         rst_controller_009_reset_out_reset;                                                                 // rst_controller_009:reset_out -> [cmd_xbar_mux_040:reset, cmd_xbar_mux_041:reset, cmd_xbar_mux_042:reset, ctod_0:reset_n, ctod_0_in_csr_translator:reset, ctod_0_in_csr_translator_avalon_universal_slave_0_agent:reset, ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ctod_0_in_translator:reset, ctod_0_in_translator_avalon_universal_slave_0_agent:reset, ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ctod_0_out_translator:reset, ctod_0_out_translator_avalon_universal_slave_0_agent:reset, ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_040:reset, id_router_041:reset, id_router_042:reset, rsp_xbar_demux_040:reset, rsp_xbar_demux_041:reset, rsp_xbar_demux_042:reset]
	wire         rst_controller_010_reset_out_reset;                                                                 // rst_controller_010:reset_out -> [cmd_xbar_mux_031:reset, cmd_xbar_mux_032:reset, cmd_xbar_mux_033:reset, dtoe_0:reset_n, dtoe_0_in_csr_translator:reset, dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:reset, dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dtoe_0_in_translator:reset, dtoe_0_in_translator_avalon_universal_slave_0_agent:reset, dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dtoe_0_out_translator:reset, dtoe_0_out_translator_avalon_universal_slave_0_agent:reset, dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_031:reset, id_router_032:reset, id_router_033:reset, rsp_xbar_demux_031:reset, rsp_xbar_demux_032:reset, rsp_xbar_demux_033:reset]
	wire         rst_controller_011_reset_out_reset;                                                                 // rst_controller_011:reset_out -> [cmd_xbar_mux_022:reset, cmd_xbar_mux_023:reset, cmd_xbar_mux_024:reset, etof_0:reset_n, etof_0_in_csr_translator:reset, etof_0_in_csr_translator_avalon_universal_slave_0_agent:reset, etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, etof_0_in_translator:reset, etof_0_in_translator_avalon_universal_slave_0_agent:reset, etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, etof_0_out_translator:reset, etof_0_out_translator_avalon_universal_slave_0_agent:reset, etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset]
	wire         rst_controller_012_reset_out_reset;                                                                 // rst_controller_012:reset_out -> [atof_0:reset_n, atof_0_in_csr_translator:reset, atof_0_in_csr_translator_avalon_universal_slave_0_agent:reset, atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atof_0_in_translator:reset, atof_0_in_translator_avalon_universal_slave_0_agent:reset, atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atof_0_out_translator:reset, atof_0_out_translator_avalon_universal_slave_0_agent:reset, atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_017:reset, cmd_xbar_mux_018:reset, cmd_xbar_mux_019:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset]
	wire         rst_controller_013_reset_out_reset;                                                                 // rst_controller_013:reset_out -> [atod_0:reset_n, atod_0_in_csr_translator:reset, atod_0_in_csr_translator_avalon_universal_slave_0_agent:reset, atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atod_0_in_translator:reset, atod_0_in_translator_avalon_universal_slave_0_agent:reset, atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atod_0_out_translator:reset, atod_0_out_translator_avalon_universal_slave_0_agent:reset, atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_011:reset, cmd_xbar_mux_012:reset, cmd_xbar_mux_013:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset]
	wire         rst_controller_014_reset_out_reset;                                                                 // rst_controller_014:reset_out -> [atoe_0:reset_n, atoe_0_in_csr_translator:reset, atoe_0_in_csr_translator_avalon_universal_slave_0_agent:reset, atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atoe_0_in_translator:reset, atoe_0_in_translator_avalon_universal_slave_0_agent:reset, atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, atoe_0_out_translator:reset, atoe_0_out_translator_avalon_universal_slave_0_agent:reset, atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_014:reset, cmd_xbar_mux_015:reset, cmd_xbar_mux_016:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                    // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                          // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                  // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src0_data;                                                                           // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [65:0] cmd_xbar_demux_src0_channel;                                                                        // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                          // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                    // cmd_xbar_demux:src1_endofpacket -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                          // cmd_xbar_demux:src1_valid -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                  // cmd_xbar_demux:src1_startofpacket -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_src1_data;                                                                           // cmd_xbar_demux:src1_data -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_src1_channel;                                                                        // cmd_xbar_demux:src1_channel -> ins_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src2_endofpacket;                                                                    // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                          // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                  // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src2_data;                                                                           // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [65:0] cmd_xbar_demux_src2_channel;                                                                        // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                          // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                    // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                          // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                  // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src3_data;                                                                           // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire  [65:0] cmd_xbar_demux_src3_channel;                                                                        // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                          // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_src4_endofpacket;                                                                    // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                          // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                  // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src4_data;                                                                           // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire  [65:0] cmd_xbar_demux_src4_channel;                                                                        // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire         cmd_xbar_demux_src4_ready;                                                                          // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire         cmd_xbar_demux_src5_endofpacket;                                                                    // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                                          // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                                  // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src5_data;                                                                           // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire  [65:0] cmd_xbar_demux_src5_channel;                                                                        // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire         cmd_xbar_demux_src5_ready;                                                                          // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire         cmd_xbar_demux_src6_endofpacket;                                                                    // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                                          // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                                  // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src6_data;                                                                           // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire  [65:0] cmd_xbar_demux_src6_channel;                                                                        // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire         cmd_xbar_demux_src6_ready;                                                                          // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire         cmd_xbar_demux_src7_endofpacket;                                                                    // cmd_xbar_demux:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire         cmd_xbar_demux_src7_valid;                                                                          // cmd_xbar_demux:src7_valid -> cmd_xbar_mux_007:sink0_valid
	wire         cmd_xbar_demux_src7_startofpacket;                                                                  // cmd_xbar_demux:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src7_data;                                                                           // cmd_xbar_demux:src7_data -> cmd_xbar_mux_007:sink0_data
	wire  [65:0] cmd_xbar_demux_src7_channel;                                                                        // cmd_xbar_demux:src7_channel -> cmd_xbar_mux_007:sink0_channel
	wire         cmd_xbar_demux_src7_ready;                                                                          // cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux:src7_ready
	wire         cmd_xbar_demux_src8_endofpacket;                                                                    // cmd_xbar_demux:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire         cmd_xbar_demux_src8_valid;                                                                          // cmd_xbar_demux:src8_valid -> cmd_xbar_mux_008:sink0_valid
	wire         cmd_xbar_demux_src8_startofpacket;                                                                  // cmd_xbar_demux:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src8_data;                                                                           // cmd_xbar_demux:src8_data -> cmd_xbar_mux_008:sink0_data
	wire  [65:0] cmd_xbar_demux_src8_channel;                                                                        // cmd_xbar_demux:src8_channel -> cmd_xbar_mux_008:sink0_channel
	wire         cmd_xbar_demux_src8_ready;                                                                          // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux:src8_ready
	wire         cmd_xbar_demux_src9_endofpacket;                                                                    // cmd_xbar_demux:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire         cmd_xbar_demux_src9_valid;                                                                          // cmd_xbar_demux:src9_valid -> cmd_xbar_mux_009:sink0_valid
	wire         cmd_xbar_demux_src9_startofpacket;                                                                  // cmd_xbar_demux:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src9_data;                                                                           // cmd_xbar_demux:src9_data -> cmd_xbar_mux_009:sink0_data
	wire  [65:0] cmd_xbar_demux_src9_channel;                                                                        // cmd_xbar_demux:src9_channel -> cmd_xbar_mux_009:sink0_channel
	wire         cmd_xbar_demux_src9_ready;                                                                          // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux:src9_ready
	wire         cmd_xbar_demux_src10_endofpacket;                                                                   // cmd_xbar_demux:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire         cmd_xbar_demux_src10_valid;                                                                         // cmd_xbar_demux:src10_valid -> cmd_xbar_mux_010:sink0_valid
	wire         cmd_xbar_demux_src10_startofpacket;                                                                 // cmd_xbar_demux:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src10_data;                                                                          // cmd_xbar_demux:src10_data -> cmd_xbar_mux_010:sink0_data
	wire  [65:0] cmd_xbar_demux_src10_channel;                                                                       // cmd_xbar_demux:src10_channel -> cmd_xbar_mux_010:sink0_channel
	wire         cmd_xbar_demux_src10_ready;                                                                         // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux:src10_ready
	wire         cmd_xbar_demux_src11_endofpacket;                                                                   // cmd_xbar_demux:src11_endofpacket -> cmd_xbar_mux_011:sink0_endofpacket
	wire         cmd_xbar_demux_src11_valid;                                                                         // cmd_xbar_demux:src11_valid -> cmd_xbar_mux_011:sink0_valid
	wire         cmd_xbar_demux_src11_startofpacket;                                                                 // cmd_xbar_demux:src11_startofpacket -> cmd_xbar_mux_011:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src11_data;                                                                          // cmd_xbar_demux:src11_data -> cmd_xbar_mux_011:sink0_data
	wire  [65:0] cmd_xbar_demux_src11_channel;                                                                       // cmd_xbar_demux:src11_channel -> cmd_xbar_mux_011:sink0_channel
	wire         cmd_xbar_demux_src11_ready;                                                                         // cmd_xbar_mux_011:sink0_ready -> cmd_xbar_demux:src11_ready
	wire         cmd_xbar_demux_src12_endofpacket;                                                                   // cmd_xbar_demux:src12_endofpacket -> cmd_xbar_mux_012:sink0_endofpacket
	wire         cmd_xbar_demux_src12_valid;                                                                         // cmd_xbar_demux:src12_valid -> cmd_xbar_mux_012:sink0_valid
	wire         cmd_xbar_demux_src12_startofpacket;                                                                 // cmd_xbar_demux:src12_startofpacket -> cmd_xbar_mux_012:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src12_data;                                                                          // cmd_xbar_demux:src12_data -> cmd_xbar_mux_012:sink0_data
	wire  [65:0] cmd_xbar_demux_src12_channel;                                                                       // cmd_xbar_demux:src12_channel -> cmd_xbar_mux_012:sink0_channel
	wire         cmd_xbar_demux_src12_ready;                                                                         // cmd_xbar_mux_012:sink0_ready -> cmd_xbar_demux:src12_ready
	wire         cmd_xbar_demux_src13_endofpacket;                                                                   // cmd_xbar_demux:src13_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	wire         cmd_xbar_demux_src13_valid;                                                                         // cmd_xbar_demux:src13_valid -> cmd_xbar_mux_013:sink0_valid
	wire         cmd_xbar_demux_src13_startofpacket;                                                                 // cmd_xbar_demux:src13_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src13_data;                                                                          // cmd_xbar_demux:src13_data -> cmd_xbar_mux_013:sink0_data
	wire  [65:0] cmd_xbar_demux_src13_channel;                                                                       // cmd_xbar_demux:src13_channel -> cmd_xbar_mux_013:sink0_channel
	wire         cmd_xbar_demux_src13_ready;                                                                         // cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux:src13_ready
	wire         cmd_xbar_demux_src14_endofpacket;                                                                   // cmd_xbar_demux:src14_endofpacket -> cmd_xbar_mux_014:sink0_endofpacket
	wire         cmd_xbar_demux_src14_valid;                                                                         // cmd_xbar_demux:src14_valid -> cmd_xbar_mux_014:sink0_valid
	wire         cmd_xbar_demux_src14_startofpacket;                                                                 // cmd_xbar_demux:src14_startofpacket -> cmd_xbar_mux_014:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src14_data;                                                                          // cmd_xbar_demux:src14_data -> cmd_xbar_mux_014:sink0_data
	wire  [65:0] cmd_xbar_demux_src14_channel;                                                                       // cmd_xbar_demux:src14_channel -> cmd_xbar_mux_014:sink0_channel
	wire         cmd_xbar_demux_src14_ready;                                                                         // cmd_xbar_mux_014:sink0_ready -> cmd_xbar_demux:src14_ready
	wire         cmd_xbar_demux_src15_endofpacket;                                                                   // cmd_xbar_demux:src15_endofpacket -> cmd_xbar_mux_015:sink0_endofpacket
	wire         cmd_xbar_demux_src15_valid;                                                                         // cmd_xbar_demux:src15_valid -> cmd_xbar_mux_015:sink0_valid
	wire         cmd_xbar_demux_src15_startofpacket;                                                                 // cmd_xbar_demux:src15_startofpacket -> cmd_xbar_mux_015:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src15_data;                                                                          // cmd_xbar_demux:src15_data -> cmd_xbar_mux_015:sink0_data
	wire  [65:0] cmd_xbar_demux_src15_channel;                                                                       // cmd_xbar_demux:src15_channel -> cmd_xbar_mux_015:sink0_channel
	wire         cmd_xbar_demux_src15_ready;                                                                         // cmd_xbar_mux_015:sink0_ready -> cmd_xbar_demux:src15_ready
	wire         cmd_xbar_demux_src16_endofpacket;                                                                   // cmd_xbar_demux:src16_endofpacket -> cmd_xbar_mux_016:sink0_endofpacket
	wire         cmd_xbar_demux_src16_valid;                                                                         // cmd_xbar_demux:src16_valid -> cmd_xbar_mux_016:sink0_valid
	wire         cmd_xbar_demux_src16_startofpacket;                                                                 // cmd_xbar_demux:src16_startofpacket -> cmd_xbar_mux_016:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src16_data;                                                                          // cmd_xbar_demux:src16_data -> cmd_xbar_mux_016:sink0_data
	wire  [65:0] cmd_xbar_demux_src16_channel;                                                                       // cmd_xbar_demux:src16_channel -> cmd_xbar_mux_016:sink0_channel
	wire         cmd_xbar_demux_src16_ready;                                                                         // cmd_xbar_mux_016:sink0_ready -> cmd_xbar_demux:src16_ready
	wire         cmd_xbar_demux_src17_endofpacket;                                                                   // cmd_xbar_demux:src17_endofpacket -> cmd_xbar_mux_017:sink0_endofpacket
	wire         cmd_xbar_demux_src17_valid;                                                                         // cmd_xbar_demux:src17_valid -> cmd_xbar_mux_017:sink0_valid
	wire         cmd_xbar_demux_src17_startofpacket;                                                                 // cmd_xbar_demux:src17_startofpacket -> cmd_xbar_mux_017:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src17_data;                                                                          // cmd_xbar_demux:src17_data -> cmd_xbar_mux_017:sink0_data
	wire  [65:0] cmd_xbar_demux_src17_channel;                                                                       // cmd_xbar_demux:src17_channel -> cmd_xbar_mux_017:sink0_channel
	wire         cmd_xbar_demux_src17_ready;                                                                         // cmd_xbar_mux_017:sink0_ready -> cmd_xbar_demux:src17_ready
	wire         cmd_xbar_demux_src18_endofpacket;                                                                   // cmd_xbar_demux:src18_endofpacket -> cmd_xbar_mux_018:sink0_endofpacket
	wire         cmd_xbar_demux_src18_valid;                                                                         // cmd_xbar_demux:src18_valid -> cmd_xbar_mux_018:sink0_valid
	wire         cmd_xbar_demux_src18_startofpacket;                                                                 // cmd_xbar_demux:src18_startofpacket -> cmd_xbar_mux_018:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src18_data;                                                                          // cmd_xbar_demux:src18_data -> cmd_xbar_mux_018:sink0_data
	wire  [65:0] cmd_xbar_demux_src18_channel;                                                                       // cmd_xbar_demux:src18_channel -> cmd_xbar_mux_018:sink0_channel
	wire         cmd_xbar_demux_src18_ready;                                                                         // cmd_xbar_mux_018:sink0_ready -> cmd_xbar_demux:src18_ready
	wire         cmd_xbar_demux_src19_endofpacket;                                                                   // cmd_xbar_demux:src19_endofpacket -> cmd_xbar_mux_019:sink0_endofpacket
	wire         cmd_xbar_demux_src19_valid;                                                                         // cmd_xbar_demux:src19_valid -> cmd_xbar_mux_019:sink0_valid
	wire         cmd_xbar_demux_src19_startofpacket;                                                                 // cmd_xbar_demux:src19_startofpacket -> cmd_xbar_mux_019:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src19_data;                                                                          // cmd_xbar_demux:src19_data -> cmd_xbar_mux_019:sink0_data
	wire  [65:0] cmd_xbar_demux_src19_channel;                                                                       // cmd_xbar_demux:src19_channel -> cmd_xbar_mux_019:sink0_channel
	wire         cmd_xbar_demux_src19_ready;                                                                         // cmd_xbar_mux_019:sink0_ready -> cmd_xbar_demux:src19_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux_017:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                      // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux_017:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                              // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux_017:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src0_data;                                                                       // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux_017:sink1_data
	wire  [65:0] cmd_xbar_demux_001_src0_channel;                                                                    // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux_017:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                      // cmd_xbar_mux_017:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_018:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                      // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_018:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                              // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_018:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src1_data;                                                                       // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_018:sink1_data
	wire  [65:0] cmd_xbar_demux_001_src1_channel;                                                                    // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_018:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                      // cmd_xbar_mux_018:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_019:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                      // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_019:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                              // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_019:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src2_data;                                                                       // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_019:sink1_data
	wire  [65:0] cmd_xbar_demux_001_src2_channel;                                                                    // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_019:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                      // cmd_xbar_mux_019:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                // cmd_xbar_demux_001:src3_endofpacket -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                      // cmd_xbar_demux_001:src3_valid -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                              // cmd_xbar_demux_001:src3_startofpacket -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src3_data;                                                                       // cmd_xbar_demux_001:src3_data -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_001_src3_channel;                                                                    // cmd_xbar_demux_001:src3_channel -> ins_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_021:sink0_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                      // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_021:sink0_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                              // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_021:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src4_data;                                                                       // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_021:sink0_data
	wire  [65:0] cmd_xbar_demux_001_src4_channel;                                                                    // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_021:sink0_channel
	wire         cmd_xbar_demux_001_src4_ready;                                                                      // cmd_xbar_mux_021:sink0_ready -> cmd_xbar_demux_001:src4_ready
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_022:sink0_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                      // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_022:sink0_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                              // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_022:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src5_data;                                                                       // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_022:sink0_data
	wire  [65:0] cmd_xbar_demux_001_src5_channel;                                                                    // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_022:sink0_channel
	wire         cmd_xbar_demux_001_src5_ready;                                                                      // cmd_xbar_mux_022:sink0_ready -> cmd_xbar_demux_001:src5_ready
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                // cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_023:sink0_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                      // cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_023:sink0_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                              // cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_023:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src6_data;                                                                       // cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_023:sink0_data
	wire  [65:0] cmd_xbar_demux_001_src6_channel;                                                                    // cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_023:sink0_channel
	wire         cmd_xbar_demux_001_src6_ready;                                                                      // cmd_xbar_mux_023:sink0_ready -> cmd_xbar_demux_001:src6_ready
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                // cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_024:sink0_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                      // cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_024:sink0_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                              // cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_024:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src7_data;                                                                       // cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_024:sink0_data
	wire  [65:0] cmd_xbar_demux_001_src7_channel;                                                                    // cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_024:sink0_channel
	wire         cmd_xbar_demux_001_src7_ready;                                                                      // cmd_xbar_mux_024:sink0_ready -> cmd_xbar_demux_001:src7_ready
	wire         cmd_xbar_demux_002_src0_endofpacket;                                                                // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_017:sink2_endofpacket
	wire         cmd_xbar_demux_002_src0_valid;                                                                      // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_017:sink2_valid
	wire         cmd_xbar_demux_002_src0_startofpacket;                                                              // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_017:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src0_data;                                                                       // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_017:sink2_data
	wire  [65:0] cmd_xbar_demux_002_src0_channel;                                                                    // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_017:sink2_channel
	wire         cmd_xbar_demux_002_src0_ready;                                                                      // cmd_xbar_mux_017:sink2_ready -> cmd_xbar_demux_002:src0_ready
	wire         cmd_xbar_demux_002_src1_endofpacket;                                                                // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_018:sink2_endofpacket
	wire         cmd_xbar_demux_002_src1_valid;                                                                      // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_018:sink2_valid
	wire         cmd_xbar_demux_002_src1_startofpacket;                                                              // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_018:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src1_data;                                                                       // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_018:sink2_data
	wire  [65:0] cmd_xbar_demux_002_src1_channel;                                                                    // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_018:sink2_channel
	wire         cmd_xbar_demux_002_src1_ready;                                                                      // cmd_xbar_mux_018:sink2_ready -> cmd_xbar_demux_002:src1_ready
	wire         cmd_xbar_demux_002_src2_endofpacket;                                                                // cmd_xbar_demux_002:src2_endofpacket -> cmd_xbar_mux_019:sink2_endofpacket
	wire         cmd_xbar_demux_002_src2_valid;                                                                      // cmd_xbar_demux_002:src2_valid -> cmd_xbar_mux_019:sink2_valid
	wire         cmd_xbar_demux_002_src2_startofpacket;                                                              // cmd_xbar_demux_002:src2_startofpacket -> cmd_xbar_mux_019:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src2_data;                                                                       // cmd_xbar_demux_002:src2_data -> cmd_xbar_mux_019:sink2_data
	wire  [65:0] cmd_xbar_demux_002_src2_channel;                                                                    // cmd_xbar_demux_002:src2_channel -> cmd_xbar_mux_019:sink2_channel
	wire         cmd_xbar_demux_002_src2_ready;                                                                      // cmd_xbar_mux_019:sink2_ready -> cmd_xbar_demux_002:src2_ready
	wire         cmd_xbar_demux_002_src3_endofpacket;                                                                // cmd_xbar_demux_002:src3_endofpacket -> cmd_xbar_mux_021:sink1_endofpacket
	wire         cmd_xbar_demux_002_src3_valid;                                                                      // cmd_xbar_demux_002:src3_valid -> cmd_xbar_mux_021:sink1_valid
	wire         cmd_xbar_demux_002_src3_startofpacket;                                                              // cmd_xbar_demux_002:src3_startofpacket -> cmd_xbar_mux_021:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src3_data;                                                                       // cmd_xbar_demux_002:src3_data -> cmd_xbar_mux_021:sink1_data
	wire  [65:0] cmd_xbar_demux_002_src3_channel;                                                                    // cmd_xbar_demux_002:src3_channel -> cmd_xbar_mux_021:sink1_channel
	wire         cmd_xbar_demux_002_src3_ready;                                                                      // cmd_xbar_mux_021:sink1_ready -> cmd_xbar_demux_002:src3_ready
	wire         cmd_xbar_demux_002_src4_endofpacket;                                                                // cmd_xbar_demux_002:src4_endofpacket -> cmd_xbar_mux_022:sink1_endofpacket
	wire         cmd_xbar_demux_002_src4_valid;                                                                      // cmd_xbar_demux_002:src4_valid -> cmd_xbar_mux_022:sink1_valid
	wire         cmd_xbar_demux_002_src4_startofpacket;                                                              // cmd_xbar_demux_002:src4_startofpacket -> cmd_xbar_mux_022:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src4_data;                                                                       // cmd_xbar_demux_002:src4_data -> cmd_xbar_mux_022:sink1_data
	wire  [65:0] cmd_xbar_demux_002_src4_channel;                                                                    // cmd_xbar_demux_002:src4_channel -> cmd_xbar_mux_022:sink1_channel
	wire         cmd_xbar_demux_002_src4_ready;                                                                      // cmd_xbar_mux_022:sink1_ready -> cmd_xbar_demux_002:src4_ready
	wire         cmd_xbar_demux_002_src5_endofpacket;                                                                // cmd_xbar_demux_002:src5_endofpacket -> cmd_xbar_mux_023:sink1_endofpacket
	wire         cmd_xbar_demux_002_src5_valid;                                                                      // cmd_xbar_demux_002:src5_valid -> cmd_xbar_mux_023:sink1_valid
	wire         cmd_xbar_demux_002_src5_startofpacket;                                                              // cmd_xbar_demux_002:src5_startofpacket -> cmd_xbar_mux_023:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src5_data;                                                                       // cmd_xbar_demux_002:src5_data -> cmd_xbar_mux_023:sink1_data
	wire  [65:0] cmd_xbar_demux_002_src5_channel;                                                                    // cmd_xbar_demux_002:src5_channel -> cmd_xbar_mux_023:sink1_channel
	wire         cmd_xbar_demux_002_src5_ready;                                                                      // cmd_xbar_mux_023:sink1_ready -> cmd_xbar_demux_002:src5_ready
	wire         cmd_xbar_demux_002_src6_endofpacket;                                                                // cmd_xbar_demux_002:src6_endofpacket -> cmd_xbar_mux_024:sink1_endofpacket
	wire         cmd_xbar_demux_002_src6_valid;                                                                      // cmd_xbar_demux_002:src6_valid -> cmd_xbar_mux_024:sink1_valid
	wire         cmd_xbar_demux_002_src6_startofpacket;                                                              // cmd_xbar_demux_002:src6_startofpacket -> cmd_xbar_mux_024:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src6_data;                                                                       // cmd_xbar_demux_002:src6_data -> cmd_xbar_mux_024:sink1_data
	wire  [65:0] cmd_xbar_demux_002_src6_channel;                                                                    // cmd_xbar_demux_002:src6_channel -> cmd_xbar_mux_024:sink1_channel
	wire         cmd_xbar_demux_002_src6_ready;                                                                      // cmd_xbar_mux_024:sink1_ready -> cmd_xbar_demux_002:src6_ready
	wire         cmd_xbar_demux_002_src7_endofpacket;                                                                // cmd_xbar_demux_002:src7_endofpacket -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src7_valid;                                                                      // cmd_xbar_demux_002:src7_valid -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src7_startofpacket;                                                              // cmd_xbar_demux_002:src7_startofpacket -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src7_data;                                                                       // cmd_xbar_demux_002:src7_data -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_002_src7_channel;                                                                    // cmd_xbar_demux_002:src7_channel -> data_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src8_endofpacket;                                                                // cmd_xbar_demux_002:src8_endofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src8_valid;                                                                      // cmd_xbar_demux_002:src8_valid -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src8_startofpacket;                                                              // cmd_xbar_demux_002:src8_startofpacket -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src8_data;                                                                       // cmd_xbar_demux_002:src8_data -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_002_src8_channel;                                                                    // cmd_xbar_demux_002:src8_channel -> jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src9_endofpacket;                                                                // cmd_xbar_demux_002:src9_endofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src9_valid;                                                                      // cmd_xbar_demux_002:src9_valid -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src9_startofpacket;                                                              // cmd_xbar_demux_002:src9_startofpacket -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src9_data;                                                                       // cmd_xbar_demux_002:src9_data -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_002_src9_channel;                                                                    // cmd_xbar_demux_002:src9_channel -> timer_5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src10_endofpacket;                                                               // cmd_xbar_demux_002:src10_endofpacket -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src10_valid;                                                                     // cmd_xbar_demux_002:src10_valid -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src10_startofpacket;                                                             // cmd_xbar_demux_002:src10_startofpacket -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_002_src10_data;                                                                      // cmd_xbar_demux_002:src10_data -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_002_src10_channel;                                                                   // cmd_xbar_demux_002:src10_channel -> high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_003_src0_endofpacket;                                                                // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_014:sink1_endofpacket
	wire         cmd_xbar_demux_003_src0_valid;                                                                      // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_014:sink1_valid
	wire         cmd_xbar_demux_003_src0_startofpacket;                                                              // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_014:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src0_data;                                                                       // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_014:sink1_data
	wire  [65:0] cmd_xbar_demux_003_src0_channel;                                                                    // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_014:sink1_channel
	wire         cmd_xbar_demux_003_src0_ready;                                                                      // cmd_xbar_mux_014:sink1_ready -> cmd_xbar_demux_003:src0_ready
	wire         cmd_xbar_demux_003_src1_endofpacket;                                                                // cmd_xbar_demux_003:src1_endofpacket -> cmd_xbar_mux_015:sink1_endofpacket
	wire         cmd_xbar_demux_003_src1_valid;                                                                      // cmd_xbar_demux_003:src1_valid -> cmd_xbar_mux_015:sink1_valid
	wire         cmd_xbar_demux_003_src1_startofpacket;                                                              // cmd_xbar_demux_003:src1_startofpacket -> cmd_xbar_mux_015:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src1_data;                                                                       // cmd_xbar_demux_003:src1_data -> cmd_xbar_mux_015:sink1_data
	wire  [65:0] cmd_xbar_demux_003_src1_channel;                                                                    // cmd_xbar_demux_003:src1_channel -> cmd_xbar_mux_015:sink1_channel
	wire         cmd_xbar_demux_003_src1_ready;                                                                      // cmd_xbar_mux_015:sink1_ready -> cmd_xbar_demux_003:src1_ready
	wire         cmd_xbar_demux_003_src2_endofpacket;                                                                // cmd_xbar_demux_003:src2_endofpacket -> cmd_xbar_mux_016:sink1_endofpacket
	wire         cmd_xbar_demux_003_src2_valid;                                                                      // cmd_xbar_demux_003:src2_valid -> cmd_xbar_mux_016:sink1_valid
	wire         cmd_xbar_demux_003_src2_startofpacket;                                                              // cmd_xbar_demux_003:src2_startofpacket -> cmd_xbar_mux_016:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src2_data;                                                                       // cmd_xbar_demux_003:src2_data -> cmd_xbar_mux_016:sink1_data
	wire  [65:0] cmd_xbar_demux_003_src2_channel;                                                                    // cmd_xbar_demux_003:src2_channel -> cmd_xbar_mux_016:sink1_channel
	wire         cmd_xbar_demux_003_src2_ready;                                                                      // cmd_xbar_mux_016:sink1_ready -> cmd_xbar_demux_003:src2_ready
	wire         cmd_xbar_demux_003_src3_endofpacket;                                                                // cmd_xbar_demux_003:src3_endofpacket -> cmd_xbar_mux_022:sink2_endofpacket
	wire         cmd_xbar_demux_003_src3_valid;                                                                      // cmd_xbar_demux_003:src3_valid -> cmd_xbar_mux_022:sink2_valid
	wire         cmd_xbar_demux_003_src3_startofpacket;                                                              // cmd_xbar_demux_003:src3_startofpacket -> cmd_xbar_mux_022:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src3_data;                                                                       // cmd_xbar_demux_003:src3_data -> cmd_xbar_mux_022:sink2_data
	wire  [65:0] cmd_xbar_demux_003_src3_channel;                                                                    // cmd_xbar_demux_003:src3_channel -> cmd_xbar_mux_022:sink2_channel
	wire         cmd_xbar_demux_003_src3_ready;                                                                      // cmd_xbar_mux_022:sink2_ready -> cmd_xbar_demux_003:src3_ready
	wire         cmd_xbar_demux_003_src4_endofpacket;                                                                // cmd_xbar_demux_003:src4_endofpacket -> cmd_xbar_mux_023:sink2_endofpacket
	wire         cmd_xbar_demux_003_src4_valid;                                                                      // cmd_xbar_demux_003:src4_valid -> cmd_xbar_mux_023:sink2_valid
	wire         cmd_xbar_demux_003_src4_startofpacket;                                                              // cmd_xbar_demux_003:src4_startofpacket -> cmd_xbar_mux_023:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src4_data;                                                                       // cmd_xbar_demux_003:src4_data -> cmd_xbar_mux_023:sink2_data
	wire  [65:0] cmd_xbar_demux_003_src4_channel;                                                                    // cmd_xbar_demux_003:src4_channel -> cmd_xbar_mux_023:sink2_channel
	wire         cmd_xbar_demux_003_src4_ready;                                                                      // cmd_xbar_mux_023:sink2_ready -> cmd_xbar_demux_003:src4_ready
	wire         cmd_xbar_demux_003_src5_endofpacket;                                                                // cmd_xbar_demux_003:src5_endofpacket -> cmd_xbar_mux_024:sink2_endofpacket
	wire         cmd_xbar_demux_003_src5_valid;                                                                      // cmd_xbar_demux_003:src5_valid -> cmd_xbar_mux_024:sink2_valid
	wire         cmd_xbar_demux_003_src5_startofpacket;                                                              // cmd_xbar_demux_003:src5_startofpacket -> cmd_xbar_mux_024:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src5_data;                                                                       // cmd_xbar_demux_003:src5_data -> cmd_xbar_mux_024:sink2_data
	wire  [65:0] cmd_xbar_demux_003_src5_channel;                                                                    // cmd_xbar_demux_003:src5_channel -> cmd_xbar_mux_024:sink2_channel
	wire         cmd_xbar_demux_003_src5_ready;                                                                      // cmd_xbar_mux_024:sink2_ready -> cmd_xbar_demux_003:src5_ready
	wire         cmd_xbar_demux_003_src6_endofpacket;                                                                // cmd_xbar_demux_003:src6_endofpacket -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_003_src6_valid;                                                                      // cmd_xbar_demux_003:src6_valid -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_003_src6_startofpacket;                                                              // cmd_xbar_demux_003:src6_startofpacket -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src6_data;                                                                       // cmd_xbar_demux_003:src6_data -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_003_src6_channel;                                                                    // cmd_xbar_demux_003:src6_channel -> ins_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_003_src7_endofpacket;                                                                // cmd_xbar_demux_003:src7_endofpacket -> cmd_xbar_mux_030:sink0_endofpacket
	wire         cmd_xbar_demux_003_src7_valid;                                                                      // cmd_xbar_demux_003:src7_valid -> cmd_xbar_mux_030:sink0_valid
	wire         cmd_xbar_demux_003_src7_startofpacket;                                                              // cmd_xbar_demux_003:src7_startofpacket -> cmd_xbar_mux_030:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src7_data;                                                                       // cmd_xbar_demux_003:src7_data -> cmd_xbar_mux_030:sink0_data
	wire  [65:0] cmd_xbar_demux_003_src7_channel;                                                                    // cmd_xbar_demux_003:src7_channel -> cmd_xbar_mux_030:sink0_channel
	wire         cmd_xbar_demux_003_src7_ready;                                                                      // cmd_xbar_mux_030:sink0_ready -> cmd_xbar_demux_003:src7_ready
	wire         cmd_xbar_demux_003_src8_endofpacket;                                                                // cmd_xbar_demux_003:src8_endofpacket -> cmd_xbar_mux_031:sink0_endofpacket
	wire         cmd_xbar_demux_003_src8_valid;                                                                      // cmd_xbar_demux_003:src8_valid -> cmd_xbar_mux_031:sink0_valid
	wire         cmd_xbar_demux_003_src8_startofpacket;                                                              // cmd_xbar_demux_003:src8_startofpacket -> cmd_xbar_mux_031:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src8_data;                                                                       // cmd_xbar_demux_003:src8_data -> cmd_xbar_mux_031:sink0_data
	wire  [65:0] cmd_xbar_demux_003_src8_channel;                                                                    // cmd_xbar_demux_003:src8_channel -> cmd_xbar_mux_031:sink0_channel
	wire         cmd_xbar_demux_003_src8_ready;                                                                      // cmd_xbar_mux_031:sink0_ready -> cmd_xbar_demux_003:src8_ready
	wire         cmd_xbar_demux_003_src9_endofpacket;                                                                // cmd_xbar_demux_003:src9_endofpacket -> cmd_xbar_mux_032:sink0_endofpacket
	wire         cmd_xbar_demux_003_src9_valid;                                                                      // cmd_xbar_demux_003:src9_valid -> cmd_xbar_mux_032:sink0_valid
	wire         cmd_xbar_demux_003_src9_startofpacket;                                                              // cmd_xbar_demux_003:src9_startofpacket -> cmd_xbar_mux_032:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src9_data;                                                                       // cmd_xbar_demux_003:src9_data -> cmd_xbar_mux_032:sink0_data
	wire  [65:0] cmd_xbar_demux_003_src9_channel;                                                                    // cmd_xbar_demux_003:src9_channel -> cmd_xbar_mux_032:sink0_channel
	wire         cmd_xbar_demux_003_src9_ready;                                                                      // cmd_xbar_mux_032:sink0_ready -> cmd_xbar_demux_003:src9_ready
	wire         cmd_xbar_demux_003_src10_endofpacket;                                                               // cmd_xbar_demux_003:src10_endofpacket -> cmd_xbar_mux_033:sink0_endofpacket
	wire         cmd_xbar_demux_003_src10_valid;                                                                     // cmd_xbar_demux_003:src10_valid -> cmd_xbar_mux_033:sink0_valid
	wire         cmd_xbar_demux_003_src10_startofpacket;                                                             // cmd_xbar_demux_003:src10_startofpacket -> cmd_xbar_mux_033:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_003_src10_data;                                                                      // cmd_xbar_demux_003:src10_data -> cmd_xbar_mux_033:sink0_data
	wire  [65:0] cmd_xbar_demux_003_src10_channel;                                                                   // cmd_xbar_demux_003:src10_channel -> cmd_xbar_mux_033:sink0_channel
	wire         cmd_xbar_demux_003_src10_ready;                                                                     // cmd_xbar_mux_033:sink0_ready -> cmd_xbar_demux_003:src10_ready
	wire         cmd_xbar_demux_004_src0_endofpacket;                                                                // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_014:sink2_endofpacket
	wire         cmd_xbar_demux_004_src0_valid;                                                                      // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_014:sink2_valid
	wire         cmd_xbar_demux_004_src0_startofpacket;                                                              // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_014:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src0_data;                                                                       // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_014:sink2_data
	wire  [65:0] cmd_xbar_demux_004_src0_channel;                                                                    // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_014:sink2_channel
	wire         cmd_xbar_demux_004_src0_ready;                                                                      // cmd_xbar_mux_014:sink2_ready -> cmd_xbar_demux_004:src0_ready
	wire         cmd_xbar_demux_004_src1_endofpacket;                                                                // cmd_xbar_demux_004:src1_endofpacket -> cmd_xbar_mux_015:sink2_endofpacket
	wire         cmd_xbar_demux_004_src1_valid;                                                                      // cmd_xbar_demux_004:src1_valid -> cmd_xbar_mux_015:sink2_valid
	wire         cmd_xbar_demux_004_src1_startofpacket;                                                              // cmd_xbar_demux_004:src1_startofpacket -> cmd_xbar_mux_015:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src1_data;                                                                       // cmd_xbar_demux_004:src1_data -> cmd_xbar_mux_015:sink2_data
	wire  [65:0] cmd_xbar_demux_004_src1_channel;                                                                    // cmd_xbar_demux_004:src1_channel -> cmd_xbar_mux_015:sink2_channel
	wire         cmd_xbar_demux_004_src1_ready;                                                                      // cmd_xbar_mux_015:sink2_ready -> cmd_xbar_demux_004:src1_ready
	wire         cmd_xbar_demux_004_src2_endofpacket;                                                                // cmd_xbar_demux_004:src2_endofpacket -> cmd_xbar_mux_016:sink2_endofpacket
	wire         cmd_xbar_demux_004_src2_valid;                                                                      // cmd_xbar_demux_004:src2_valid -> cmd_xbar_mux_016:sink2_valid
	wire         cmd_xbar_demux_004_src2_startofpacket;                                                              // cmd_xbar_demux_004:src2_startofpacket -> cmd_xbar_mux_016:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src2_data;                                                                       // cmd_xbar_demux_004:src2_data -> cmd_xbar_mux_016:sink2_data
	wire  [65:0] cmd_xbar_demux_004_src2_channel;                                                                    // cmd_xbar_demux_004:src2_channel -> cmd_xbar_mux_016:sink2_channel
	wire         cmd_xbar_demux_004_src2_ready;                                                                      // cmd_xbar_mux_016:sink2_ready -> cmd_xbar_demux_004:src2_ready
	wire         cmd_xbar_demux_004_src3_endofpacket;                                                                // cmd_xbar_demux_004:src3_endofpacket -> cmd_xbar_mux_022:sink3_endofpacket
	wire         cmd_xbar_demux_004_src3_valid;                                                                      // cmd_xbar_demux_004:src3_valid -> cmd_xbar_mux_022:sink3_valid
	wire         cmd_xbar_demux_004_src3_startofpacket;                                                              // cmd_xbar_demux_004:src3_startofpacket -> cmd_xbar_mux_022:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src3_data;                                                                       // cmd_xbar_demux_004:src3_data -> cmd_xbar_mux_022:sink3_data
	wire  [65:0] cmd_xbar_demux_004_src3_channel;                                                                    // cmd_xbar_demux_004:src3_channel -> cmd_xbar_mux_022:sink3_channel
	wire         cmd_xbar_demux_004_src3_ready;                                                                      // cmd_xbar_mux_022:sink3_ready -> cmd_xbar_demux_004:src3_ready
	wire         cmd_xbar_demux_004_src4_endofpacket;                                                                // cmd_xbar_demux_004:src4_endofpacket -> cmd_xbar_mux_023:sink3_endofpacket
	wire         cmd_xbar_demux_004_src4_valid;                                                                      // cmd_xbar_demux_004:src4_valid -> cmd_xbar_mux_023:sink3_valid
	wire         cmd_xbar_demux_004_src4_startofpacket;                                                              // cmd_xbar_demux_004:src4_startofpacket -> cmd_xbar_mux_023:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src4_data;                                                                       // cmd_xbar_demux_004:src4_data -> cmd_xbar_mux_023:sink3_data
	wire  [65:0] cmd_xbar_demux_004_src4_channel;                                                                    // cmd_xbar_demux_004:src4_channel -> cmd_xbar_mux_023:sink3_channel
	wire         cmd_xbar_demux_004_src4_ready;                                                                      // cmd_xbar_mux_023:sink3_ready -> cmd_xbar_demux_004:src4_ready
	wire         cmd_xbar_demux_004_src5_endofpacket;                                                                // cmd_xbar_demux_004:src5_endofpacket -> cmd_xbar_mux_024:sink3_endofpacket
	wire         cmd_xbar_demux_004_src5_valid;                                                                      // cmd_xbar_demux_004:src5_valid -> cmd_xbar_mux_024:sink3_valid
	wire         cmd_xbar_demux_004_src5_startofpacket;                                                              // cmd_xbar_demux_004:src5_startofpacket -> cmd_xbar_mux_024:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src5_data;                                                                       // cmd_xbar_demux_004:src5_data -> cmd_xbar_mux_024:sink3_data
	wire  [65:0] cmd_xbar_demux_004_src5_channel;                                                                    // cmd_xbar_demux_004:src5_channel -> cmd_xbar_mux_024:sink3_channel
	wire         cmd_xbar_demux_004_src5_ready;                                                                      // cmd_xbar_mux_024:sink3_ready -> cmd_xbar_demux_004:src5_ready
	wire         cmd_xbar_demux_004_src6_endofpacket;                                                                // cmd_xbar_demux_004:src6_endofpacket -> cmd_xbar_mux_030:sink1_endofpacket
	wire         cmd_xbar_demux_004_src6_valid;                                                                      // cmd_xbar_demux_004:src6_valid -> cmd_xbar_mux_030:sink1_valid
	wire         cmd_xbar_demux_004_src6_startofpacket;                                                              // cmd_xbar_demux_004:src6_startofpacket -> cmd_xbar_mux_030:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src6_data;                                                                       // cmd_xbar_demux_004:src6_data -> cmd_xbar_mux_030:sink1_data
	wire  [65:0] cmd_xbar_demux_004_src6_channel;                                                                    // cmd_xbar_demux_004:src6_channel -> cmd_xbar_mux_030:sink1_channel
	wire         cmd_xbar_demux_004_src6_ready;                                                                      // cmd_xbar_mux_030:sink1_ready -> cmd_xbar_demux_004:src6_ready
	wire         cmd_xbar_demux_004_src7_endofpacket;                                                                // cmd_xbar_demux_004:src7_endofpacket -> cmd_xbar_mux_031:sink1_endofpacket
	wire         cmd_xbar_demux_004_src7_valid;                                                                      // cmd_xbar_demux_004:src7_valid -> cmd_xbar_mux_031:sink1_valid
	wire         cmd_xbar_demux_004_src7_startofpacket;                                                              // cmd_xbar_demux_004:src7_startofpacket -> cmd_xbar_mux_031:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src7_data;                                                                       // cmd_xbar_demux_004:src7_data -> cmd_xbar_mux_031:sink1_data
	wire  [65:0] cmd_xbar_demux_004_src7_channel;                                                                    // cmd_xbar_demux_004:src7_channel -> cmd_xbar_mux_031:sink1_channel
	wire         cmd_xbar_demux_004_src7_ready;                                                                      // cmd_xbar_mux_031:sink1_ready -> cmd_xbar_demux_004:src7_ready
	wire         cmd_xbar_demux_004_src8_endofpacket;                                                                // cmd_xbar_demux_004:src8_endofpacket -> cmd_xbar_mux_032:sink1_endofpacket
	wire         cmd_xbar_demux_004_src8_valid;                                                                      // cmd_xbar_demux_004:src8_valid -> cmd_xbar_mux_032:sink1_valid
	wire         cmd_xbar_demux_004_src8_startofpacket;                                                              // cmd_xbar_demux_004:src8_startofpacket -> cmd_xbar_mux_032:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src8_data;                                                                       // cmd_xbar_demux_004:src8_data -> cmd_xbar_mux_032:sink1_data
	wire  [65:0] cmd_xbar_demux_004_src8_channel;                                                                    // cmd_xbar_demux_004:src8_channel -> cmd_xbar_mux_032:sink1_channel
	wire         cmd_xbar_demux_004_src8_ready;                                                                      // cmd_xbar_mux_032:sink1_ready -> cmd_xbar_demux_004:src8_ready
	wire         cmd_xbar_demux_004_src9_endofpacket;                                                                // cmd_xbar_demux_004:src9_endofpacket -> cmd_xbar_mux_033:sink1_endofpacket
	wire         cmd_xbar_demux_004_src9_valid;                                                                      // cmd_xbar_demux_004:src9_valid -> cmd_xbar_mux_033:sink1_valid
	wire         cmd_xbar_demux_004_src9_startofpacket;                                                              // cmd_xbar_demux_004:src9_startofpacket -> cmd_xbar_mux_033:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src9_data;                                                                       // cmd_xbar_demux_004:src9_data -> cmd_xbar_mux_033:sink1_data
	wire  [65:0] cmd_xbar_demux_004_src9_channel;                                                                    // cmd_xbar_demux_004:src9_channel -> cmd_xbar_mux_033:sink1_channel
	wire         cmd_xbar_demux_004_src9_ready;                                                                      // cmd_xbar_mux_033:sink1_ready -> cmd_xbar_demux_004:src9_ready
	wire         cmd_xbar_demux_004_src10_endofpacket;                                                               // cmd_xbar_demux_004:src10_endofpacket -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src10_valid;                                                                     // cmd_xbar_demux_004:src10_valid -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src10_startofpacket;                                                             // cmd_xbar_demux_004:src10_startofpacket -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src10_data;                                                                      // cmd_xbar_demux_004:src10_data -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_004_src10_channel;                                                                   // cmd_xbar_demux_004:src10_channel -> data_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src11_endofpacket;                                                               // cmd_xbar_demux_004:src11_endofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src11_valid;                                                                     // cmd_xbar_demux_004:src11_valid -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src11_startofpacket;                                                             // cmd_xbar_demux_004:src11_startofpacket -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src11_data;                                                                      // cmd_xbar_demux_004:src11_data -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_004_src11_channel;                                                                   // cmd_xbar_demux_004:src11_channel -> jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src12_endofpacket;                                                               // cmd_xbar_demux_004:src12_endofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src12_valid;                                                                     // cmd_xbar_demux_004:src12_valid -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src12_startofpacket;                                                             // cmd_xbar_demux_004:src12_startofpacket -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src12_data;                                                                      // cmd_xbar_demux_004:src12_data -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_004_src12_channel;                                                                   // cmd_xbar_demux_004:src12_channel -> timer_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src13_endofpacket;                                                               // cmd_xbar_demux_004:src13_endofpacket -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src13_valid;                                                                     // cmd_xbar_demux_004:src13_valid -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src13_startofpacket;                                                             // cmd_xbar_demux_004:src13_startofpacket -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_004_src13_data;                                                                      // cmd_xbar_demux_004:src13_data -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_004_src13_channel;                                                                   // cmd_xbar_demux_004:src13_channel -> high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_005_src0_endofpacket;                                                                // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_011:sink1_endofpacket
	wire         cmd_xbar_demux_005_src0_valid;                                                                      // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_011:sink1_valid
	wire         cmd_xbar_demux_005_src0_startofpacket;                                                              // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_011:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src0_data;                                                                       // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_011:sink1_data
	wire  [65:0] cmd_xbar_demux_005_src0_channel;                                                                    // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_011:sink1_channel
	wire         cmd_xbar_demux_005_src0_ready;                                                                      // cmd_xbar_mux_011:sink1_ready -> cmd_xbar_demux_005:src0_ready
	wire         cmd_xbar_demux_005_src1_endofpacket;                                                                // cmd_xbar_demux_005:src1_endofpacket -> cmd_xbar_mux_012:sink1_endofpacket
	wire         cmd_xbar_demux_005_src1_valid;                                                                      // cmd_xbar_demux_005:src1_valid -> cmd_xbar_mux_012:sink1_valid
	wire         cmd_xbar_demux_005_src1_startofpacket;                                                              // cmd_xbar_demux_005:src1_startofpacket -> cmd_xbar_mux_012:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src1_data;                                                                       // cmd_xbar_demux_005:src1_data -> cmd_xbar_mux_012:sink1_data
	wire  [65:0] cmd_xbar_demux_005_src1_channel;                                                                    // cmd_xbar_demux_005:src1_channel -> cmd_xbar_mux_012:sink1_channel
	wire         cmd_xbar_demux_005_src1_ready;                                                                      // cmd_xbar_mux_012:sink1_ready -> cmd_xbar_demux_005:src1_ready
	wire         cmd_xbar_demux_005_src2_endofpacket;                                                                // cmd_xbar_demux_005:src2_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	wire         cmd_xbar_demux_005_src2_valid;                                                                      // cmd_xbar_demux_005:src2_valid -> cmd_xbar_mux_013:sink1_valid
	wire         cmd_xbar_demux_005_src2_startofpacket;                                                              // cmd_xbar_demux_005:src2_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src2_data;                                                                       // cmd_xbar_demux_005:src2_data -> cmd_xbar_mux_013:sink1_data
	wire  [65:0] cmd_xbar_demux_005_src2_channel;                                                                    // cmd_xbar_demux_005:src2_channel -> cmd_xbar_mux_013:sink1_channel
	wire         cmd_xbar_demux_005_src2_ready;                                                                      // cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_005:src2_ready
	wire         cmd_xbar_demux_005_src3_endofpacket;                                                                // cmd_xbar_demux_005:src3_endofpacket -> cmd_xbar_mux_031:sink2_endofpacket
	wire         cmd_xbar_demux_005_src3_valid;                                                                      // cmd_xbar_demux_005:src3_valid -> cmd_xbar_mux_031:sink2_valid
	wire         cmd_xbar_demux_005_src3_startofpacket;                                                              // cmd_xbar_demux_005:src3_startofpacket -> cmd_xbar_mux_031:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src3_data;                                                                       // cmd_xbar_demux_005:src3_data -> cmd_xbar_mux_031:sink2_data
	wire  [65:0] cmd_xbar_demux_005_src3_channel;                                                                    // cmd_xbar_demux_005:src3_channel -> cmd_xbar_mux_031:sink2_channel
	wire         cmd_xbar_demux_005_src3_ready;                                                                      // cmd_xbar_mux_031:sink2_ready -> cmd_xbar_demux_005:src3_ready
	wire         cmd_xbar_demux_005_src4_endofpacket;                                                                // cmd_xbar_demux_005:src4_endofpacket -> cmd_xbar_mux_032:sink2_endofpacket
	wire         cmd_xbar_demux_005_src4_valid;                                                                      // cmd_xbar_demux_005:src4_valid -> cmd_xbar_mux_032:sink2_valid
	wire         cmd_xbar_demux_005_src4_startofpacket;                                                              // cmd_xbar_demux_005:src4_startofpacket -> cmd_xbar_mux_032:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src4_data;                                                                       // cmd_xbar_demux_005:src4_data -> cmd_xbar_mux_032:sink2_data
	wire  [65:0] cmd_xbar_demux_005_src4_channel;                                                                    // cmd_xbar_demux_005:src4_channel -> cmd_xbar_mux_032:sink2_channel
	wire         cmd_xbar_demux_005_src4_ready;                                                                      // cmd_xbar_mux_032:sink2_ready -> cmd_xbar_demux_005:src4_ready
	wire         cmd_xbar_demux_005_src5_endofpacket;                                                                // cmd_xbar_demux_005:src5_endofpacket -> cmd_xbar_mux_033:sink2_endofpacket
	wire         cmd_xbar_demux_005_src5_valid;                                                                      // cmd_xbar_demux_005:src5_valid -> cmd_xbar_mux_033:sink2_valid
	wire         cmd_xbar_demux_005_src5_startofpacket;                                                              // cmd_xbar_demux_005:src5_startofpacket -> cmd_xbar_mux_033:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src5_data;                                                                       // cmd_xbar_demux_005:src5_data -> cmd_xbar_mux_033:sink2_data
	wire  [65:0] cmd_xbar_demux_005_src5_channel;                                                                    // cmd_xbar_demux_005:src5_channel -> cmd_xbar_mux_033:sink2_channel
	wire         cmd_xbar_demux_005_src5_ready;                                                                      // cmd_xbar_mux_033:sink2_ready -> cmd_xbar_demux_005:src5_ready
	wire         cmd_xbar_demux_005_src6_endofpacket;                                                                // cmd_xbar_demux_005:src6_endofpacket -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_005_src6_valid;                                                                      // cmd_xbar_demux_005:src6_valid -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_005_src6_startofpacket;                                                              // cmd_xbar_demux_005:src6_startofpacket -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src6_data;                                                                       // cmd_xbar_demux_005:src6_data -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_005_src6_channel;                                                                    // cmd_xbar_demux_005:src6_channel -> ins_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_005_src7_endofpacket;                                                                // cmd_xbar_demux_005:src7_endofpacket -> cmd_xbar_mux_039:sink0_endofpacket
	wire         cmd_xbar_demux_005_src7_valid;                                                                      // cmd_xbar_demux_005:src7_valid -> cmd_xbar_mux_039:sink0_valid
	wire         cmd_xbar_demux_005_src7_startofpacket;                                                              // cmd_xbar_demux_005:src7_startofpacket -> cmd_xbar_mux_039:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src7_data;                                                                       // cmd_xbar_demux_005:src7_data -> cmd_xbar_mux_039:sink0_data
	wire  [65:0] cmd_xbar_demux_005_src7_channel;                                                                    // cmd_xbar_demux_005:src7_channel -> cmd_xbar_mux_039:sink0_channel
	wire         cmd_xbar_demux_005_src7_ready;                                                                      // cmd_xbar_mux_039:sink0_ready -> cmd_xbar_demux_005:src7_ready
	wire         cmd_xbar_demux_005_src8_endofpacket;                                                                // cmd_xbar_demux_005:src8_endofpacket -> cmd_xbar_mux_040:sink0_endofpacket
	wire         cmd_xbar_demux_005_src8_valid;                                                                      // cmd_xbar_demux_005:src8_valid -> cmd_xbar_mux_040:sink0_valid
	wire         cmd_xbar_demux_005_src8_startofpacket;                                                              // cmd_xbar_demux_005:src8_startofpacket -> cmd_xbar_mux_040:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src8_data;                                                                       // cmd_xbar_demux_005:src8_data -> cmd_xbar_mux_040:sink0_data
	wire  [65:0] cmd_xbar_demux_005_src8_channel;                                                                    // cmd_xbar_demux_005:src8_channel -> cmd_xbar_mux_040:sink0_channel
	wire         cmd_xbar_demux_005_src8_ready;                                                                      // cmd_xbar_mux_040:sink0_ready -> cmd_xbar_demux_005:src8_ready
	wire         cmd_xbar_demux_005_src9_endofpacket;                                                                // cmd_xbar_demux_005:src9_endofpacket -> cmd_xbar_mux_041:sink0_endofpacket
	wire         cmd_xbar_demux_005_src9_valid;                                                                      // cmd_xbar_demux_005:src9_valid -> cmd_xbar_mux_041:sink0_valid
	wire         cmd_xbar_demux_005_src9_startofpacket;                                                              // cmd_xbar_demux_005:src9_startofpacket -> cmd_xbar_mux_041:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src9_data;                                                                       // cmd_xbar_demux_005:src9_data -> cmd_xbar_mux_041:sink0_data
	wire  [65:0] cmd_xbar_demux_005_src9_channel;                                                                    // cmd_xbar_demux_005:src9_channel -> cmd_xbar_mux_041:sink0_channel
	wire         cmd_xbar_demux_005_src9_ready;                                                                      // cmd_xbar_mux_041:sink0_ready -> cmd_xbar_demux_005:src9_ready
	wire         cmd_xbar_demux_005_src10_endofpacket;                                                               // cmd_xbar_demux_005:src10_endofpacket -> cmd_xbar_mux_042:sink0_endofpacket
	wire         cmd_xbar_demux_005_src10_valid;                                                                     // cmd_xbar_demux_005:src10_valid -> cmd_xbar_mux_042:sink0_valid
	wire         cmd_xbar_demux_005_src10_startofpacket;                                                             // cmd_xbar_demux_005:src10_startofpacket -> cmd_xbar_mux_042:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_005_src10_data;                                                                      // cmd_xbar_demux_005:src10_data -> cmd_xbar_mux_042:sink0_data
	wire  [65:0] cmd_xbar_demux_005_src10_channel;                                                                   // cmd_xbar_demux_005:src10_channel -> cmd_xbar_mux_042:sink0_channel
	wire         cmd_xbar_demux_005_src10_ready;                                                                     // cmd_xbar_mux_042:sink0_ready -> cmd_xbar_demux_005:src10_ready
	wire         cmd_xbar_demux_006_src0_endofpacket;                                                                // cmd_xbar_demux_006:src0_endofpacket -> cmd_xbar_mux_011:sink2_endofpacket
	wire         cmd_xbar_demux_006_src0_valid;                                                                      // cmd_xbar_demux_006:src0_valid -> cmd_xbar_mux_011:sink2_valid
	wire         cmd_xbar_demux_006_src0_startofpacket;                                                              // cmd_xbar_demux_006:src0_startofpacket -> cmd_xbar_mux_011:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src0_data;                                                                       // cmd_xbar_demux_006:src0_data -> cmd_xbar_mux_011:sink2_data
	wire  [65:0] cmd_xbar_demux_006_src0_channel;                                                                    // cmd_xbar_demux_006:src0_channel -> cmd_xbar_mux_011:sink2_channel
	wire         cmd_xbar_demux_006_src0_ready;                                                                      // cmd_xbar_mux_011:sink2_ready -> cmd_xbar_demux_006:src0_ready
	wire         cmd_xbar_demux_006_src1_endofpacket;                                                                // cmd_xbar_demux_006:src1_endofpacket -> cmd_xbar_mux_012:sink2_endofpacket
	wire         cmd_xbar_demux_006_src1_valid;                                                                      // cmd_xbar_demux_006:src1_valid -> cmd_xbar_mux_012:sink2_valid
	wire         cmd_xbar_demux_006_src1_startofpacket;                                                              // cmd_xbar_demux_006:src1_startofpacket -> cmd_xbar_mux_012:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src1_data;                                                                       // cmd_xbar_demux_006:src1_data -> cmd_xbar_mux_012:sink2_data
	wire  [65:0] cmd_xbar_demux_006_src1_channel;                                                                    // cmd_xbar_demux_006:src1_channel -> cmd_xbar_mux_012:sink2_channel
	wire         cmd_xbar_demux_006_src1_ready;                                                                      // cmd_xbar_mux_012:sink2_ready -> cmd_xbar_demux_006:src1_ready
	wire         cmd_xbar_demux_006_src2_endofpacket;                                                                // cmd_xbar_demux_006:src2_endofpacket -> cmd_xbar_mux_013:sink2_endofpacket
	wire         cmd_xbar_demux_006_src2_valid;                                                                      // cmd_xbar_demux_006:src2_valid -> cmd_xbar_mux_013:sink2_valid
	wire         cmd_xbar_demux_006_src2_startofpacket;                                                              // cmd_xbar_demux_006:src2_startofpacket -> cmd_xbar_mux_013:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src2_data;                                                                       // cmd_xbar_demux_006:src2_data -> cmd_xbar_mux_013:sink2_data
	wire  [65:0] cmd_xbar_demux_006_src2_channel;                                                                    // cmd_xbar_demux_006:src2_channel -> cmd_xbar_mux_013:sink2_channel
	wire         cmd_xbar_demux_006_src2_ready;                                                                      // cmd_xbar_mux_013:sink2_ready -> cmd_xbar_demux_006:src2_ready
	wire         cmd_xbar_demux_006_src3_endofpacket;                                                                // cmd_xbar_demux_006:src3_endofpacket -> cmd_xbar_mux_031:sink3_endofpacket
	wire         cmd_xbar_demux_006_src3_valid;                                                                      // cmd_xbar_demux_006:src3_valid -> cmd_xbar_mux_031:sink3_valid
	wire         cmd_xbar_demux_006_src3_startofpacket;                                                              // cmd_xbar_demux_006:src3_startofpacket -> cmd_xbar_mux_031:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src3_data;                                                                       // cmd_xbar_demux_006:src3_data -> cmd_xbar_mux_031:sink3_data
	wire  [65:0] cmd_xbar_demux_006_src3_channel;                                                                    // cmd_xbar_demux_006:src3_channel -> cmd_xbar_mux_031:sink3_channel
	wire         cmd_xbar_demux_006_src3_ready;                                                                      // cmd_xbar_mux_031:sink3_ready -> cmd_xbar_demux_006:src3_ready
	wire         cmd_xbar_demux_006_src4_endofpacket;                                                                // cmd_xbar_demux_006:src4_endofpacket -> cmd_xbar_mux_032:sink3_endofpacket
	wire         cmd_xbar_demux_006_src4_valid;                                                                      // cmd_xbar_demux_006:src4_valid -> cmd_xbar_mux_032:sink3_valid
	wire         cmd_xbar_demux_006_src4_startofpacket;                                                              // cmd_xbar_demux_006:src4_startofpacket -> cmd_xbar_mux_032:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src4_data;                                                                       // cmd_xbar_demux_006:src4_data -> cmd_xbar_mux_032:sink3_data
	wire  [65:0] cmd_xbar_demux_006_src4_channel;                                                                    // cmd_xbar_demux_006:src4_channel -> cmd_xbar_mux_032:sink3_channel
	wire         cmd_xbar_demux_006_src4_ready;                                                                      // cmd_xbar_mux_032:sink3_ready -> cmd_xbar_demux_006:src4_ready
	wire         cmd_xbar_demux_006_src5_endofpacket;                                                                // cmd_xbar_demux_006:src5_endofpacket -> cmd_xbar_mux_033:sink3_endofpacket
	wire         cmd_xbar_demux_006_src5_valid;                                                                      // cmd_xbar_demux_006:src5_valid -> cmd_xbar_mux_033:sink3_valid
	wire         cmd_xbar_demux_006_src5_startofpacket;                                                              // cmd_xbar_demux_006:src5_startofpacket -> cmd_xbar_mux_033:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src5_data;                                                                       // cmd_xbar_demux_006:src5_data -> cmd_xbar_mux_033:sink3_data
	wire  [65:0] cmd_xbar_demux_006_src5_channel;                                                                    // cmd_xbar_demux_006:src5_channel -> cmd_xbar_mux_033:sink3_channel
	wire         cmd_xbar_demux_006_src5_ready;                                                                      // cmd_xbar_mux_033:sink3_ready -> cmd_xbar_demux_006:src5_ready
	wire         cmd_xbar_demux_006_src6_endofpacket;                                                                // cmd_xbar_demux_006:src6_endofpacket -> cmd_xbar_mux_039:sink1_endofpacket
	wire         cmd_xbar_demux_006_src6_valid;                                                                      // cmd_xbar_demux_006:src6_valid -> cmd_xbar_mux_039:sink1_valid
	wire         cmd_xbar_demux_006_src6_startofpacket;                                                              // cmd_xbar_demux_006:src6_startofpacket -> cmd_xbar_mux_039:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src6_data;                                                                       // cmd_xbar_demux_006:src6_data -> cmd_xbar_mux_039:sink1_data
	wire  [65:0] cmd_xbar_demux_006_src6_channel;                                                                    // cmd_xbar_demux_006:src6_channel -> cmd_xbar_mux_039:sink1_channel
	wire         cmd_xbar_demux_006_src6_ready;                                                                      // cmd_xbar_mux_039:sink1_ready -> cmd_xbar_demux_006:src6_ready
	wire         cmd_xbar_demux_006_src7_endofpacket;                                                                // cmd_xbar_demux_006:src7_endofpacket -> cmd_xbar_mux_040:sink1_endofpacket
	wire         cmd_xbar_demux_006_src7_valid;                                                                      // cmd_xbar_demux_006:src7_valid -> cmd_xbar_mux_040:sink1_valid
	wire         cmd_xbar_demux_006_src7_startofpacket;                                                              // cmd_xbar_demux_006:src7_startofpacket -> cmd_xbar_mux_040:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src7_data;                                                                       // cmd_xbar_demux_006:src7_data -> cmd_xbar_mux_040:sink1_data
	wire  [65:0] cmd_xbar_demux_006_src7_channel;                                                                    // cmd_xbar_demux_006:src7_channel -> cmd_xbar_mux_040:sink1_channel
	wire         cmd_xbar_demux_006_src7_ready;                                                                      // cmd_xbar_mux_040:sink1_ready -> cmd_xbar_demux_006:src7_ready
	wire         cmd_xbar_demux_006_src8_endofpacket;                                                                // cmd_xbar_demux_006:src8_endofpacket -> cmd_xbar_mux_041:sink1_endofpacket
	wire         cmd_xbar_demux_006_src8_valid;                                                                      // cmd_xbar_demux_006:src8_valid -> cmd_xbar_mux_041:sink1_valid
	wire         cmd_xbar_demux_006_src8_startofpacket;                                                              // cmd_xbar_demux_006:src8_startofpacket -> cmd_xbar_mux_041:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src8_data;                                                                       // cmd_xbar_demux_006:src8_data -> cmd_xbar_mux_041:sink1_data
	wire  [65:0] cmd_xbar_demux_006_src8_channel;                                                                    // cmd_xbar_demux_006:src8_channel -> cmd_xbar_mux_041:sink1_channel
	wire         cmd_xbar_demux_006_src8_ready;                                                                      // cmd_xbar_mux_041:sink1_ready -> cmd_xbar_demux_006:src8_ready
	wire         cmd_xbar_demux_006_src9_endofpacket;                                                                // cmd_xbar_demux_006:src9_endofpacket -> cmd_xbar_mux_042:sink1_endofpacket
	wire         cmd_xbar_demux_006_src9_valid;                                                                      // cmd_xbar_demux_006:src9_valid -> cmd_xbar_mux_042:sink1_valid
	wire         cmd_xbar_demux_006_src9_startofpacket;                                                              // cmd_xbar_demux_006:src9_startofpacket -> cmd_xbar_mux_042:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src9_data;                                                                       // cmd_xbar_demux_006:src9_data -> cmd_xbar_mux_042:sink1_data
	wire  [65:0] cmd_xbar_demux_006_src9_channel;                                                                    // cmd_xbar_demux_006:src9_channel -> cmd_xbar_mux_042:sink1_channel
	wire         cmd_xbar_demux_006_src9_ready;                                                                      // cmd_xbar_mux_042:sink1_ready -> cmd_xbar_demux_006:src9_ready
	wire         cmd_xbar_demux_006_src10_endofpacket;                                                               // cmd_xbar_demux_006:src10_endofpacket -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_006_src10_valid;                                                                     // cmd_xbar_demux_006:src10_valid -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_006_src10_startofpacket;                                                             // cmd_xbar_demux_006:src10_startofpacket -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src10_data;                                                                      // cmd_xbar_demux_006:src10_data -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_006_src10_channel;                                                                   // cmd_xbar_demux_006:src10_channel -> data_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_006_src11_endofpacket;                                                               // cmd_xbar_demux_006:src11_endofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_006_src11_valid;                                                                     // cmd_xbar_demux_006:src11_valid -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_006_src11_startofpacket;                                                             // cmd_xbar_demux_006:src11_startofpacket -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src11_data;                                                                      // cmd_xbar_demux_006:src11_data -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_006_src11_channel;                                                                   // cmd_xbar_demux_006:src11_channel -> jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_006_src12_endofpacket;                                                               // cmd_xbar_demux_006:src12_endofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_006_src12_valid;                                                                     // cmd_xbar_demux_006:src12_valid -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_006_src12_startofpacket;                                                             // cmd_xbar_demux_006:src12_startofpacket -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src12_data;                                                                      // cmd_xbar_demux_006:src12_data -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_006_src12_channel;                                                                   // cmd_xbar_demux_006:src12_channel -> timer_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_006_src13_endofpacket;                                                               // cmd_xbar_demux_006:src13_endofpacket -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_006_src13_valid;                                                                     // cmd_xbar_demux_006:src13_valid -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_006_src13_startofpacket;                                                             // cmd_xbar_demux_006:src13_startofpacket -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_006_src13_data;                                                                      // cmd_xbar_demux_006:src13_data -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_006_src13_channel;                                                                   // cmd_xbar_demux_006:src13_channel -> high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_007_src0_endofpacket;                                                                // cmd_xbar_demux_007:src0_endofpacket -> cmd_xbar_mux_040:sink2_endofpacket
	wire         cmd_xbar_demux_007_src0_valid;                                                                      // cmd_xbar_demux_007:src0_valid -> cmd_xbar_mux_040:sink2_valid
	wire         cmd_xbar_demux_007_src0_startofpacket;                                                              // cmd_xbar_demux_007:src0_startofpacket -> cmd_xbar_mux_040:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src0_data;                                                                       // cmd_xbar_demux_007:src0_data -> cmd_xbar_mux_040:sink2_data
	wire  [65:0] cmd_xbar_demux_007_src0_channel;                                                                    // cmd_xbar_demux_007:src0_channel -> cmd_xbar_mux_040:sink2_channel
	wire         cmd_xbar_demux_007_src0_ready;                                                                      // cmd_xbar_mux_040:sink2_ready -> cmd_xbar_demux_007:src0_ready
	wire         cmd_xbar_demux_007_src1_endofpacket;                                                                // cmd_xbar_demux_007:src1_endofpacket -> cmd_xbar_mux_041:sink2_endofpacket
	wire         cmd_xbar_demux_007_src1_valid;                                                                      // cmd_xbar_demux_007:src1_valid -> cmd_xbar_mux_041:sink2_valid
	wire         cmd_xbar_demux_007_src1_startofpacket;                                                              // cmd_xbar_demux_007:src1_startofpacket -> cmd_xbar_mux_041:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src1_data;                                                                       // cmd_xbar_demux_007:src1_data -> cmd_xbar_mux_041:sink2_data
	wire  [65:0] cmd_xbar_demux_007_src1_channel;                                                                    // cmd_xbar_demux_007:src1_channel -> cmd_xbar_mux_041:sink2_channel
	wire         cmd_xbar_demux_007_src1_ready;                                                                      // cmd_xbar_mux_041:sink2_ready -> cmd_xbar_demux_007:src1_ready
	wire         cmd_xbar_demux_007_src2_endofpacket;                                                                // cmd_xbar_demux_007:src2_endofpacket -> cmd_xbar_mux_042:sink2_endofpacket
	wire         cmd_xbar_demux_007_src2_valid;                                                                      // cmd_xbar_demux_007:src2_valid -> cmd_xbar_mux_042:sink2_valid
	wire         cmd_xbar_demux_007_src2_startofpacket;                                                              // cmd_xbar_demux_007:src2_startofpacket -> cmd_xbar_mux_042:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src2_data;                                                                       // cmd_xbar_demux_007:src2_data -> cmd_xbar_mux_042:sink2_data
	wire  [65:0] cmd_xbar_demux_007_src2_channel;                                                                    // cmd_xbar_demux_007:src2_channel -> cmd_xbar_mux_042:sink2_channel
	wire         cmd_xbar_demux_007_src2_ready;                                                                      // cmd_xbar_mux_042:sink2_ready -> cmd_xbar_demux_007:src2_ready
	wire         cmd_xbar_demux_007_src3_endofpacket;                                                                // cmd_xbar_demux_007:src3_endofpacket -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_007_src3_valid;                                                                      // cmd_xbar_demux_007:src3_valid -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_007_src3_startofpacket;                                                              // cmd_xbar_demux_007:src3_startofpacket -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src3_data;                                                                       // cmd_xbar_demux_007:src3_data -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_007_src3_channel;                                                                    // cmd_xbar_demux_007:src3_channel -> data_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_007_src4_endofpacket;                                                                // cmd_xbar_demux_007:src4_endofpacket -> cmd_xbar_mux_048:sink0_endofpacket
	wire         cmd_xbar_demux_007_src4_valid;                                                                      // cmd_xbar_demux_007:src4_valid -> cmd_xbar_mux_048:sink0_valid
	wire         cmd_xbar_demux_007_src4_startofpacket;                                                              // cmd_xbar_demux_007:src4_startofpacket -> cmd_xbar_mux_048:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src4_data;                                                                       // cmd_xbar_demux_007:src4_data -> cmd_xbar_mux_048:sink0_data
	wire  [65:0] cmd_xbar_demux_007_src4_channel;                                                                    // cmd_xbar_demux_007:src4_channel -> cmd_xbar_mux_048:sink0_channel
	wire         cmd_xbar_demux_007_src4_ready;                                                                      // cmd_xbar_mux_048:sink0_ready -> cmd_xbar_demux_007:src4_ready
	wire         cmd_xbar_demux_007_src5_endofpacket;                                                                // cmd_xbar_demux_007:src5_endofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_007_src5_valid;                                                                      // cmd_xbar_demux_007:src5_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_007_src5_startofpacket;                                                              // cmd_xbar_demux_007:src5_startofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src5_data;                                                                       // cmd_xbar_demux_007:src5_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_007_src5_channel;                                                                    // cmd_xbar_demux_007:src5_channel -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_007_src6_endofpacket;                                                                // cmd_xbar_demux_007:src6_endofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_007_src6_valid;                                                                      // cmd_xbar_demux_007:src6_valid -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_007_src6_startofpacket;                                                              // cmd_xbar_demux_007:src6_startofpacket -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src6_data;                                                                       // cmd_xbar_demux_007:src6_data -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_007_src6_channel;                                                                    // cmd_xbar_demux_007:src6_channel -> timer_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_007_src7_endofpacket;                                                                // cmd_xbar_demux_007:src7_endofpacket -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_007_src7_valid;                                                                      // cmd_xbar_demux_007:src7_valid -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_007_src7_startofpacket;                                                              // cmd_xbar_demux_007:src7_startofpacket -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src7_data;                                                                       // cmd_xbar_demux_007:src7_data -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_007_src7_channel;                                                                    // cmd_xbar_demux_007:src7_channel -> high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_007_src8_endofpacket;                                                                // cmd_xbar_demux_007:src8_endofpacket -> cmd_xbar_mux_052:sink0_endofpacket
	wire         cmd_xbar_demux_007_src8_valid;                                                                      // cmd_xbar_demux_007:src8_valid -> cmd_xbar_mux_052:sink0_valid
	wire         cmd_xbar_demux_007_src8_startofpacket;                                                              // cmd_xbar_demux_007:src8_startofpacket -> cmd_xbar_mux_052:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src8_data;                                                                       // cmd_xbar_demux_007:src8_data -> cmd_xbar_mux_052:sink0_data
	wire  [65:0] cmd_xbar_demux_007_src8_channel;                                                                    // cmd_xbar_demux_007:src8_channel -> cmd_xbar_mux_052:sink0_channel
	wire         cmd_xbar_demux_007_src8_ready;                                                                      // cmd_xbar_mux_052:sink0_ready -> cmd_xbar_demux_007:src8_ready
	wire         cmd_xbar_demux_007_src9_endofpacket;                                                                // cmd_xbar_demux_007:src9_endofpacket -> cmd_xbar_mux_053:sink0_endofpacket
	wire         cmd_xbar_demux_007_src9_valid;                                                                      // cmd_xbar_demux_007:src9_valid -> cmd_xbar_mux_053:sink0_valid
	wire         cmd_xbar_demux_007_src9_startofpacket;                                                              // cmd_xbar_demux_007:src9_startofpacket -> cmd_xbar_mux_053:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src9_data;                                                                       // cmd_xbar_demux_007:src9_data -> cmd_xbar_mux_053:sink0_data
	wire  [65:0] cmd_xbar_demux_007_src9_channel;                                                                    // cmd_xbar_demux_007:src9_channel -> cmd_xbar_mux_053:sink0_channel
	wire         cmd_xbar_demux_007_src9_ready;                                                                      // cmd_xbar_mux_053:sink0_ready -> cmd_xbar_demux_007:src9_ready
	wire         cmd_xbar_demux_007_src10_endofpacket;                                                               // cmd_xbar_demux_007:src10_endofpacket -> cmd_xbar_mux_054:sink0_endofpacket
	wire         cmd_xbar_demux_007_src10_valid;                                                                     // cmd_xbar_demux_007:src10_valid -> cmd_xbar_mux_054:sink0_valid
	wire         cmd_xbar_demux_007_src10_startofpacket;                                                             // cmd_xbar_demux_007:src10_startofpacket -> cmd_xbar_mux_054:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_007_src10_data;                                                                      // cmd_xbar_demux_007:src10_data -> cmd_xbar_mux_054:sink0_data
	wire  [65:0] cmd_xbar_demux_007_src10_channel;                                                                   // cmd_xbar_demux_007:src10_channel -> cmd_xbar_mux_054:sink0_channel
	wire         cmd_xbar_demux_007_src10_ready;                                                                     // cmd_xbar_mux_054:sink0_ready -> cmd_xbar_demux_007:src10_ready
	wire         cmd_xbar_demux_008_src0_endofpacket;                                                                // cmd_xbar_demux_008:src0_endofpacket -> cmd_xbar_mux_040:sink3_endofpacket
	wire         cmd_xbar_demux_008_src0_valid;                                                                      // cmd_xbar_demux_008:src0_valid -> cmd_xbar_mux_040:sink3_valid
	wire         cmd_xbar_demux_008_src0_startofpacket;                                                              // cmd_xbar_demux_008:src0_startofpacket -> cmd_xbar_mux_040:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_008_src0_data;                                                                       // cmd_xbar_demux_008:src0_data -> cmd_xbar_mux_040:sink3_data
	wire  [65:0] cmd_xbar_demux_008_src0_channel;                                                                    // cmd_xbar_demux_008:src0_channel -> cmd_xbar_mux_040:sink3_channel
	wire         cmd_xbar_demux_008_src0_ready;                                                                      // cmd_xbar_mux_040:sink3_ready -> cmd_xbar_demux_008:src0_ready
	wire         cmd_xbar_demux_008_src1_endofpacket;                                                                // cmd_xbar_demux_008:src1_endofpacket -> cmd_xbar_mux_041:sink3_endofpacket
	wire         cmd_xbar_demux_008_src1_valid;                                                                      // cmd_xbar_demux_008:src1_valid -> cmd_xbar_mux_041:sink3_valid
	wire         cmd_xbar_demux_008_src1_startofpacket;                                                              // cmd_xbar_demux_008:src1_startofpacket -> cmd_xbar_mux_041:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_008_src1_data;                                                                       // cmd_xbar_demux_008:src1_data -> cmd_xbar_mux_041:sink3_data
	wire  [65:0] cmd_xbar_demux_008_src1_channel;                                                                    // cmd_xbar_demux_008:src1_channel -> cmd_xbar_mux_041:sink3_channel
	wire         cmd_xbar_demux_008_src1_ready;                                                                      // cmd_xbar_mux_041:sink3_ready -> cmd_xbar_demux_008:src1_ready
	wire         cmd_xbar_demux_008_src2_endofpacket;                                                                // cmd_xbar_demux_008:src2_endofpacket -> cmd_xbar_mux_042:sink3_endofpacket
	wire         cmd_xbar_demux_008_src2_valid;                                                                      // cmd_xbar_demux_008:src2_valid -> cmd_xbar_mux_042:sink3_valid
	wire         cmd_xbar_demux_008_src2_startofpacket;                                                              // cmd_xbar_demux_008:src2_startofpacket -> cmd_xbar_mux_042:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_008_src2_data;                                                                       // cmd_xbar_demux_008:src2_data -> cmd_xbar_mux_042:sink3_data
	wire  [65:0] cmd_xbar_demux_008_src2_channel;                                                                    // cmd_xbar_demux_008:src2_channel -> cmd_xbar_mux_042:sink3_channel
	wire         cmd_xbar_demux_008_src2_ready;                                                                      // cmd_xbar_mux_042:sink3_ready -> cmd_xbar_demux_008:src2_ready
	wire         cmd_xbar_demux_008_src3_endofpacket;                                                                // cmd_xbar_demux_008:src3_endofpacket -> cmd_xbar_mux_048:sink1_endofpacket
	wire         cmd_xbar_demux_008_src3_valid;                                                                      // cmd_xbar_demux_008:src3_valid -> cmd_xbar_mux_048:sink1_valid
	wire         cmd_xbar_demux_008_src3_startofpacket;                                                              // cmd_xbar_demux_008:src3_startofpacket -> cmd_xbar_mux_048:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_008_src3_data;                                                                       // cmd_xbar_demux_008:src3_data -> cmd_xbar_mux_048:sink1_data
	wire  [65:0] cmd_xbar_demux_008_src3_channel;                                                                    // cmd_xbar_demux_008:src3_channel -> cmd_xbar_mux_048:sink1_channel
	wire         cmd_xbar_demux_008_src3_ready;                                                                      // cmd_xbar_mux_048:sink1_ready -> cmd_xbar_demux_008:src3_ready
	wire         cmd_xbar_demux_008_src4_endofpacket;                                                                // cmd_xbar_demux_008:src4_endofpacket -> cmd_xbar_mux_052:sink1_endofpacket
	wire         cmd_xbar_demux_008_src4_valid;                                                                      // cmd_xbar_demux_008:src4_valid -> cmd_xbar_mux_052:sink1_valid
	wire         cmd_xbar_demux_008_src4_startofpacket;                                                              // cmd_xbar_demux_008:src4_startofpacket -> cmd_xbar_mux_052:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_008_src4_data;                                                                       // cmd_xbar_demux_008:src4_data -> cmd_xbar_mux_052:sink1_data
	wire  [65:0] cmd_xbar_demux_008_src4_channel;                                                                    // cmd_xbar_demux_008:src4_channel -> cmd_xbar_mux_052:sink1_channel
	wire         cmd_xbar_demux_008_src4_ready;                                                                      // cmd_xbar_mux_052:sink1_ready -> cmd_xbar_demux_008:src4_ready
	wire         cmd_xbar_demux_008_src5_endofpacket;                                                                // cmd_xbar_demux_008:src5_endofpacket -> cmd_xbar_mux_053:sink1_endofpacket
	wire         cmd_xbar_demux_008_src5_valid;                                                                      // cmd_xbar_demux_008:src5_valid -> cmd_xbar_mux_053:sink1_valid
	wire         cmd_xbar_demux_008_src5_startofpacket;                                                              // cmd_xbar_demux_008:src5_startofpacket -> cmd_xbar_mux_053:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_008_src5_data;                                                                       // cmd_xbar_demux_008:src5_data -> cmd_xbar_mux_053:sink1_data
	wire  [65:0] cmd_xbar_demux_008_src5_channel;                                                                    // cmd_xbar_demux_008:src5_channel -> cmd_xbar_mux_053:sink1_channel
	wire         cmd_xbar_demux_008_src5_ready;                                                                      // cmd_xbar_mux_053:sink1_ready -> cmd_xbar_demux_008:src5_ready
	wire         cmd_xbar_demux_008_src6_endofpacket;                                                                // cmd_xbar_demux_008:src6_endofpacket -> cmd_xbar_mux_054:sink1_endofpacket
	wire         cmd_xbar_demux_008_src6_valid;                                                                      // cmd_xbar_demux_008:src6_valid -> cmd_xbar_mux_054:sink1_valid
	wire         cmd_xbar_demux_008_src6_startofpacket;                                                              // cmd_xbar_demux_008:src6_startofpacket -> cmd_xbar_mux_054:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_008_src6_data;                                                                       // cmd_xbar_demux_008:src6_data -> cmd_xbar_mux_054:sink1_data
	wire  [65:0] cmd_xbar_demux_008_src6_channel;                                                                    // cmd_xbar_demux_008:src6_channel -> cmd_xbar_mux_054:sink1_channel
	wire         cmd_xbar_demux_008_src6_ready;                                                                      // cmd_xbar_mux_054:sink1_ready -> cmd_xbar_demux_008:src6_ready
	wire         cmd_xbar_demux_008_src7_endofpacket;                                                                // cmd_xbar_demux_008:src7_endofpacket -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_008_src7_valid;                                                                      // cmd_xbar_demux_008:src7_valid -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_008_src7_startofpacket;                                                              // cmd_xbar_demux_008:src7_startofpacket -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_008_src7_data;                                                                       // cmd_xbar_demux_008:src7_data -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_008_src7_channel;                                                                    // cmd_xbar_demux_008:src7_channel -> ins_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_009_src0_endofpacket;                                                                // cmd_xbar_demux_009:src0_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_009_src0_valid;                                                                      // cmd_xbar_demux_009:src0_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_009_src0_startofpacket;                                                              // cmd_xbar_demux_009:src0_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src0_data;                                                                       // cmd_xbar_demux_009:src0_data -> cmd_xbar_mux_002:sink1_data
	wire  [65:0] cmd_xbar_demux_009_src0_channel;                                                                    // cmd_xbar_demux_009:src0_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_009_src0_ready;                                                                      // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_009:src0_ready
	wire         cmd_xbar_demux_009_src1_endofpacket;                                                                // cmd_xbar_demux_009:src1_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_009_src1_valid;                                                                      // cmd_xbar_demux_009:src1_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_009_src1_startofpacket;                                                              // cmd_xbar_demux_009:src1_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src1_data;                                                                       // cmd_xbar_demux_009:src1_data -> cmd_xbar_mux_003:sink1_data
	wire  [65:0] cmd_xbar_demux_009_src1_channel;                                                                    // cmd_xbar_demux_009:src1_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_009_src1_ready;                                                                      // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_009:src1_ready
	wire         cmd_xbar_demux_009_src2_endofpacket;                                                                // cmd_xbar_demux_009:src2_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire         cmd_xbar_demux_009_src2_valid;                                                                      // cmd_xbar_demux_009:src2_valid -> cmd_xbar_mux_004:sink1_valid
	wire         cmd_xbar_demux_009_src2_startofpacket;                                                              // cmd_xbar_demux_009:src2_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src2_data;                                                                       // cmd_xbar_demux_009:src2_data -> cmd_xbar_mux_004:sink1_data
	wire  [65:0] cmd_xbar_demux_009_src2_channel;                                                                    // cmd_xbar_demux_009:src2_channel -> cmd_xbar_mux_004:sink1_channel
	wire         cmd_xbar_demux_009_src2_ready;                                                                      // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_009:src2_ready
	wire         cmd_xbar_demux_009_src3_endofpacket;                                                                // cmd_xbar_demux_009:src3_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire         cmd_xbar_demux_009_src3_valid;                                                                      // cmd_xbar_demux_009:src3_valid -> cmd_xbar_mux_005:sink1_valid
	wire         cmd_xbar_demux_009_src3_startofpacket;                                                              // cmd_xbar_demux_009:src3_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src3_data;                                                                       // cmd_xbar_demux_009:src3_data -> cmd_xbar_mux_005:sink1_data
	wire  [65:0] cmd_xbar_demux_009_src3_channel;                                                                    // cmd_xbar_demux_009:src3_channel -> cmd_xbar_mux_005:sink1_channel
	wire         cmd_xbar_demux_009_src3_ready;                                                                      // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_009:src3_ready
	wire         cmd_xbar_demux_009_src4_endofpacket;                                                                // cmd_xbar_demux_009:src4_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire         cmd_xbar_demux_009_src4_valid;                                                                      // cmd_xbar_demux_009:src4_valid -> cmd_xbar_mux_006:sink1_valid
	wire         cmd_xbar_demux_009_src4_startofpacket;                                                              // cmd_xbar_demux_009:src4_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src4_data;                                                                       // cmd_xbar_demux_009:src4_data -> cmd_xbar_mux_006:sink1_data
	wire  [65:0] cmd_xbar_demux_009_src4_channel;                                                                    // cmd_xbar_demux_009:src4_channel -> cmd_xbar_mux_006:sink1_channel
	wire         cmd_xbar_demux_009_src4_ready;                                                                      // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_009:src4_ready
	wire         cmd_xbar_demux_009_src5_endofpacket;                                                                // cmd_xbar_demux_009:src5_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire         cmd_xbar_demux_009_src5_valid;                                                                      // cmd_xbar_demux_009:src5_valid -> cmd_xbar_mux_007:sink1_valid
	wire         cmd_xbar_demux_009_src5_startofpacket;                                                              // cmd_xbar_demux_009:src5_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src5_data;                                                                       // cmd_xbar_demux_009:src5_data -> cmd_xbar_mux_007:sink1_data
	wire  [65:0] cmd_xbar_demux_009_src5_channel;                                                                    // cmd_xbar_demux_009:src5_channel -> cmd_xbar_mux_007:sink1_channel
	wire         cmd_xbar_demux_009_src5_ready;                                                                      // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_009:src5_ready
	wire         cmd_xbar_demux_009_src6_endofpacket;                                                                // cmd_xbar_demux_009:src6_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire         cmd_xbar_demux_009_src6_valid;                                                                      // cmd_xbar_demux_009:src6_valid -> cmd_xbar_mux_008:sink1_valid
	wire         cmd_xbar_demux_009_src6_startofpacket;                                                              // cmd_xbar_demux_009:src6_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src6_data;                                                                       // cmd_xbar_demux_009:src6_data -> cmd_xbar_mux_008:sink1_data
	wire  [65:0] cmd_xbar_demux_009_src6_channel;                                                                    // cmd_xbar_demux_009:src6_channel -> cmd_xbar_mux_008:sink1_channel
	wire         cmd_xbar_demux_009_src6_ready;                                                                      // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_009:src6_ready
	wire         cmd_xbar_demux_009_src7_endofpacket;                                                                // cmd_xbar_demux_009:src7_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire         cmd_xbar_demux_009_src7_valid;                                                                      // cmd_xbar_demux_009:src7_valid -> cmd_xbar_mux_009:sink1_valid
	wire         cmd_xbar_demux_009_src7_startofpacket;                                                              // cmd_xbar_demux_009:src7_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src7_data;                                                                       // cmd_xbar_demux_009:src7_data -> cmd_xbar_mux_009:sink1_data
	wire  [65:0] cmd_xbar_demux_009_src7_channel;                                                                    // cmd_xbar_demux_009:src7_channel -> cmd_xbar_mux_009:sink1_channel
	wire         cmd_xbar_demux_009_src7_ready;                                                                      // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_009:src7_ready
	wire         cmd_xbar_demux_009_src8_endofpacket;                                                                // cmd_xbar_demux_009:src8_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire         cmd_xbar_demux_009_src8_valid;                                                                      // cmd_xbar_demux_009:src8_valid -> cmd_xbar_mux_010:sink1_valid
	wire         cmd_xbar_demux_009_src8_startofpacket;                                                              // cmd_xbar_demux_009:src8_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src8_data;                                                                       // cmd_xbar_demux_009:src8_data -> cmd_xbar_mux_010:sink1_data
	wire  [65:0] cmd_xbar_demux_009_src8_channel;                                                                    // cmd_xbar_demux_009:src8_channel -> cmd_xbar_mux_010:sink1_channel
	wire         cmd_xbar_demux_009_src8_ready;                                                                      // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_009:src8_ready
	wire         cmd_xbar_demux_009_src9_endofpacket;                                                                // cmd_xbar_demux_009:src9_endofpacket -> cmd_xbar_mux_052:sink2_endofpacket
	wire         cmd_xbar_demux_009_src9_valid;                                                                      // cmd_xbar_demux_009:src9_valid -> cmd_xbar_mux_052:sink2_valid
	wire         cmd_xbar_demux_009_src9_startofpacket;                                                              // cmd_xbar_demux_009:src9_startofpacket -> cmd_xbar_mux_052:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src9_data;                                                                       // cmd_xbar_demux_009:src9_data -> cmd_xbar_mux_052:sink2_data
	wire  [65:0] cmd_xbar_demux_009_src9_channel;                                                                    // cmd_xbar_demux_009:src9_channel -> cmd_xbar_mux_052:sink2_channel
	wire         cmd_xbar_demux_009_src9_ready;                                                                      // cmd_xbar_mux_052:sink2_ready -> cmd_xbar_demux_009:src9_ready
	wire         cmd_xbar_demux_009_src10_endofpacket;                                                               // cmd_xbar_demux_009:src10_endofpacket -> cmd_xbar_mux_053:sink2_endofpacket
	wire         cmd_xbar_demux_009_src10_valid;                                                                     // cmd_xbar_demux_009:src10_valid -> cmd_xbar_mux_053:sink2_valid
	wire         cmd_xbar_demux_009_src10_startofpacket;                                                             // cmd_xbar_demux_009:src10_startofpacket -> cmd_xbar_mux_053:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src10_data;                                                                      // cmd_xbar_demux_009:src10_data -> cmd_xbar_mux_053:sink2_data
	wire  [65:0] cmd_xbar_demux_009_src10_channel;                                                                   // cmd_xbar_demux_009:src10_channel -> cmd_xbar_mux_053:sink2_channel
	wire         cmd_xbar_demux_009_src10_ready;                                                                     // cmd_xbar_mux_053:sink2_ready -> cmd_xbar_demux_009:src10_ready
	wire         cmd_xbar_demux_009_src11_endofpacket;                                                               // cmd_xbar_demux_009:src11_endofpacket -> cmd_xbar_mux_054:sink2_endofpacket
	wire         cmd_xbar_demux_009_src11_valid;                                                                     // cmd_xbar_demux_009:src11_valid -> cmd_xbar_mux_054:sink2_valid
	wire         cmd_xbar_demux_009_src11_startofpacket;                                                             // cmd_xbar_demux_009:src11_startofpacket -> cmd_xbar_mux_054:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src11_data;                                                                      // cmd_xbar_demux_009:src11_data -> cmd_xbar_mux_054:sink2_data
	wire  [65:0] cmd_xbar_demux_009_src11_channel;                                                                   // cmd_xbar_demux_009:src11_channel -> cmd_xbar_mux_054:sink2_channel
	wire         cmd_xbar_demux_009_src11_ready;                                                                     // cmd_xbar_mux_054:sink2_ready -> cmd_xbar_demux_009:src11_ready
	wire         cmd_xbar_demux_009_src12_endofpacket;                                                               // cmd_xbar_demux_009:src12_endofpacket -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_009_src12_valid;                                                                     // cmd_xbar_demux_009:src12_valid -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_009_src12_startofpacket;                                                             // cmd_xbar_demux_009:src12_startofpacket -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src12_data;                                                                      // cmd_xbar_demux_009:src12_data -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_009_src12_channel;                                                                   // cmd_xbar_demux_009:src12_channel -> ins_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_009_src13_endofpacket;                                                               // cmd_xbar_demux_009:src13_endofpacket -> cmd_xbar_mux_057:sink0_endofpacket
	wire         cmd_xbar_demux_009_src13_valid;                                                                     // cmd_xbar_demux_009:src13_valid -> cmd_xbar_mux_057:sink0_valid
	wire         cmd_xbar_demux_009_src13_startofpacket;                                                             // cmd_xbar_demux_009:src13_startofpacket -> cmd_xbar_mux_057:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_009_src13_data;                                                                      // cmd_xbar_demux_009:src13_data -> cmd_xbar_mux_057:sink0_data
	wire  [65:0] cmd_xbar_demux_009_src13_channel;                                                                   // cmd_xbar_demux_009:src13_channel -> cmd_xbar_mux_057:sink0_channel
	wire         cmd_xbar_demux_009_src13_ready;                                                                     // cmd_xbar_mux_057:sink0_ready -> cmd_xbar_demux_009:src13_ready
	wire         cmd_xbar_demux_010_src0_endofpacket;                                                                // cmd_xbar_demux_010:src0_endofpacket -> cmd_xbar_mux_002:sink2_endofpacket
	wire         cmd_xbar_demux_010_src0_valid;                                                                      // cmd_xbar_demux_010:src0_valid -> cmd_xbar_mux_002:sink2_valid
	wire         cmd_xbar_demux_010_src0_startofpacket;                                                              // cmd_xbar_demux_010:src0_startofpacket -> cmd_xbar_mux_002:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src0_data;                                                                       // cmd_xbar_demux_010:src0_data -> cmd_xbar_mux_002:sink2_data
	wire  [65:0] cmd_xbar_demux_010_src0_channel;                                                                    // cmd_xbar_demux_010:src0_channel -> cmd_xbar_mux_002:sink2_channel
	wire         cmd_xbar_demux_010_src0_ready;                                                                      // cmd_xbar_mux_002:sink2_ready -> cmd_xbar_demux_010:src0_ready
	wire         cmd_xbar_demux_010_src1_endofpacket;                                                                // cmd_xbar_demux_010:src1_endofpacket -> cmd_xbar_mux_003:sink2_endofpacket
	wire         cmd_xbar_demux_010_src1_valid;                                                                      // cmd_xbar_demux_010:src1_valid -> cmd_xbar_mux_003:sink2_valid
	wire         cmd_xbar_demux_010_src1_startofpacket;                                                              // cmd_xbar_demux_010:src1_startofpacket -> cmd_xbar_mux_003:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src1_data;                                                                       // cmd_xbar_demux_010:src1_data -> cmd_xbar_mux_003:sink2_data
	wire  [65:0] cmd_xbar_demux_010_src1_channel;                                                                    // cmd_xbar_demux_010:src1_channel -> cmd_xbar_mux_003:sink2_channel
	wire         cmd_xbar_demux_010_src1_ready;                                                                      // cmd_xbar_mux_003:sink2_ready -> cmd_xbar_demux_010:src1_ready
	wire         cmd_xbar_demux_010_src2_endofpacket;                                                                // cmd_xbar_demux_010:src2_endofpacket -> cmd_xbar_mux_004:sink2_endofpacket
	wire         cmd_xbar_demux_010_src2_valid;                                                                      // cmd_xbar_demux_010:src2_valid -> cmd_xbar_mux_004:sink2_valid
	wire         cmd_xbar_demux_010_src2_startofpacket;                                                              // cmd_xbar_demux_010:src2_startofpacket -> cmd_xbar_mux_004:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src2_data;                                                                       // cmd_xbar_demux_010:src2_data -> cmd_xbar_mux_004:sink2_data
	wire  [65:0] cmd_xbar_demux_010_src2_channel;                                                                    // cmd_xbar_demux_010:src2_channel -> cmd_xbar_mux_004:sink2_channel
	wire         cmd_xbar_demux_010_src2_ready;                                                                      // cmd_xbar_mux_004:sink2_ready -> cmd_xbar_demux_010:src2_ready
	wire         cmd_xbar_demux_010_src3_endofpacket;                                                                // cmd_xbar_demux_010:src3_endofpacket -> cmd_xbar_mux_005:sink2_endofpacket
	wire         cmd_xbar_demux_010_src3_valid;                                                                      // cmd_xbar_demux_010:src3_valid -> cmd_xbar_mux_005:sink2_valid
	wire         cmd_xbar_demux_010_src3_startofpacket;                                                              // cmd_xbar_demux_010:src3_startofpacket -> cmd_xbar_mux_005:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src3_data;                                                                       // cmd_xbar_demux_010:src3_data -> cmd_xbar_mux_005:sink2_data
	wire  [65:0] cmd_xbar_demux_010_src3_channel;                                                                    // cmd_xbar_demux_010:src3_channel -> cmd_xbar_mux_005:sink2_channel
	wire         cmd_xbar_demux_010_src3_ready;                                                                      // cmd_xbar_mux_005:sink2_ready -> cmd_xbar_demux_010:src3_ready
	wire         cmd_xbar_demux_010_src4_endofpacket;                                                                // cmd_xbar_demux_010:src4_endofpacket -> cmd_xbar_mux_006:sink2_endofpacket
	wire         cmd_xbar_demux_010_src4_valid;                                                                      // cmd_xbar_demux_010:src4_valid -> cmd_xbar_mux_006:sink2_valid
	wire         cmd_xbar_demux_010_src4_startofpacket;                                                              // cmd_xbar_demux_010:src4_startofpacket -> cmd_xbar_mux_006:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src4_data;                                                                       // cmd_xbar_demux_010:src4_data -> cmd_xbar_mux_006:sink2_data
	wire  [65:0] cmd_xbar_demux_010_src4_channel;                                                                    // cmd_xbar_demux_010:src4_channel -> cmd_xbar_mux_006:sink2_channel
	wire         cmd_xbar_demux_010_src4_ready;                                                                      // cmd_xbar_mux_006:sink2_ready -> cmd_xbar_demux_010:src4_ready
	wire         cmd_xbar_demux_010_src5_endofpacket;                                                                // cmd_xbar_demux_010:src5_endofpacket -> cmd_xbar_mux_007:sink2_endofpacket
	wire         cmd_xbar_demux_010_src5_valid;                                                                      // cmd_xbar_demux_010:src5_valid -> cmd_xbar_mux_007:sink2_valid
	wire         cmd_xbar_demux_010_src5_startofpacket;                                                              // cmd_xbar_demux_010:src5_startofpacket -> cmd_xbar_mux_007:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src5_data;                                                                       // cmd_xbar_demux_010:src5_data -> cmd_xbar_mux_007:sink2_data
	wire  [65:0] cmd_xbar_demux_010_src5_channel;                                                                    // cmd_xbar_demux_010:src5_channel -> cmd_xbar_mux_007:sink2_channel
	wire         cmd_xbar_demux_010_src5_ready;                                                                      // cmd_xbar_mux_007:sink2_ready -> cmd_xbar_demux_010:src5_ready
	wire         cmd_xbar_demux_010_src6_endofpacket;                                                                // cmd_xbar_demux_010:src6_endofpacket -> cmd_xbar_mux_008:sink2_endofpacket
	wire         cmd_xbar_demux_010_src6_valid;                                                                      // cmd_xbar_demux_010:src6_valid -> cmd_xbar_mux_008:sink2_valid
	wire         cmd_xbar_demux_010_src6_startofpacket;                                                              // cmd_xbar_demux_010:src6_startofpacket -> cmd_xbar_mux_008:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src6_data;                                                                       // cmd_xbar_demux_010:src6_data -> cmd_xbar_mux_008:sink2_data
	wire  [65:0] cmd_xbar_demux_010_src6_channel;                                                                    // cmd_xbar_demux_010:src6_channel -> cmd_xbar_mux_008:sink2_channel
	wire         cmd_xbar_demux_010_src6_ready;                                                                      // cmd_xbar_mux_008:sink2_ready -> cmd_xbar_demux_010:src6_ready
	wire         cmd_xbar_demux_010_src7_endofpacket;                                                                // cmd_xbar_demux_010:src7_endofpacket -> cmd_xbar_mux_009:sink2_endofpacket
	wire         cmd_xbar_demux_010_src7_valid;                                                                      // cmd_xbar_demux_010:src7_valid -> cmd_xbar_mux_009:sink2_valid
	wire         cmd_xbar_demux_010_src7_startofpacket;                                                              // cmd_xbar_demux_010:src7_startofpacket -> cmd_xbar_mux_009:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src7_data;                                                                       // cmd_xbar_demux_010:src7_data -> cmd_xbar_mux_009:sink2_data
	wire  [65:0] cmd_xbar_demux_010_src7_channel;                                                                    // cmd_xbar_demux_010:src7_channel -> cmd_xbar_mux_009:sink2_channel
	wire         cmd_xbar_demux_010_src7_ready;                                                                      // cmd_xbar_mux_009:sink2_ready -> cmd_xbar_demux_010:src7_ready
	wire         cmd_xbar_demux_010_src8_endofpacket;                                                                // cmd_xbar_demux_010:src8_endofpacket -> cmd_xbar_mux_010:sink2_endofpacket
	wire         cmd_xbar_demux_010_src8_valid;                                                                      // cmd_xbar_demux_010:src8_valid -> cmd_xbar_mux_010:sink2_valid
	wire         cmd_xbar_demux_010_src8_startofpacket;                                                              // cmd_xbar_demux_010:src8_startofpacket -> cmd_xbar_mux_010:sink2_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src8_data;                                                                       // cmd_xbar_demux_010:src8_data -> cmd_xbar_mux_010:sink2_data
	wire  [65:0] cmd_xbar_demux_010_src8_channel;                                                                    // cmd_xbar_demux_010:src8_channel -> cmd_xbar_mux_010:sink2_channel
	wire         cmd_xbar_demux_010_src8_ready;                                                                      // cmd_xbar_mux_010:sink2_ready -> cmd_xbar_demux_010:src8_ready
	wire         cmd_xbar_demux_010_src9_endofpacket;                                                                // cmd_xbar_demux_010:src9_endofpacket -> cmd_xbar_mux_052:sink3_endofpacket
	wire         cmd_xbar_demux_010_src9_valid;                                                                      // cmd_xbar_demux_010:src9_valid -> cmd_xbar_mux_052:sink3_valid
	wire         cmd_xbar_demux_010_src9_startofpacket;                                                              // cmd_xbar_demux_010:src9_startofpacket -> cmd_xbar_mux_052:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src9_data;                                                                       // cmd_xbar_demux_010:src9_data -> cmd_xbar_mux_052:sink3_data
	wire  [65:0] cmd_xbar_demux_010_src9_channel;                                                                    // cmd_xbar_demux_010:src9_channel -> cmd_xbar_mux_052:sink3_channel
	wire         cmd_xbar_demux_010_src9_ready;                                                                      // cmd_xbar_mux_052:sink3_ready -> cmd_xbar_demux_010:src9_ready
	wire         cmd_xbar_demux_010_src10_endofpacket;                                                               // cmd_xbar_demux_010:src10_endofpacket -> cmd_xbar_mux_053:sink3_endofpacket
	wire         cmd_xbar_demux_010_src10_valid;                                                                     // cmd_xbar_demux_010:src10_valid -> cmd_xbar_mux_053:sink3_valid
	wire         cmd_xbar_demux_010_src10_startofpacket;                                                             // cmd_xbar_demux_010:src10_startofpacket -> cmd_xbar_mux_053:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src10_data;                                                                      // cmd_xbar_demux_010:src10_data -> cmd_xbar_mux_053:sink3_data
	wire  [65:0] cmd_xbar_demux_010_src10_channel;                                                                   // cmd_xbar_demux_010:src10_channel -> cmd_xbar_mux_053:sink3_channel
	wire         cmd_xbar_demux_010_src10_ready;                                                                     // cmd_xbar_mux_053:sink3_ready -> cmd_xbar_demux_010:src10_ready
	wire         cmd_xbar_demux_010_src11_endofpacket;                                                               // cmd_xbar_demux_010:src11_endofpacket -> cmd_xbar_mux_054:sink3_endofpacket
	wire         cmd_xbar_demux_010_src11_valid;                                                                     // cmd_xbar_demux_010:src11_valid -> cmd_xbar_mux_054:sink3_valid
	wire         cmd_xbar_demux_010_src11_startofpacket;                                                             // cmd_xbar_demux_010:src11_startofpacket -> cmd_xbar_mux_054:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src11_data;                                                                      // cmd_xbar_demux_010:src11_data -> cmd_xbar_mux_054:sink3_data
	wire  [65:0] cmd_xbar_demux_010_src11_channel;                                                                   // cmd_xbar_demux_010:src11_channel -> cmd_xbar_mux_054:sink3_channel
	wire         cmd_xbar_demux_010_src11_ready;                                                                     // cmd_xbar_mux_054:sink3_ready -> cmd_xbar_demux_010:src11_ready
	wire         cmd_xbar_demux_010_src12_endofpacket;                                                               // cmd_xbar_demux_010:src12_endofpacket -> cmd_xbar_mux_057:sink1_endofpacket
	wire         cmd_xbar_demux_010_src12_valid;                                                                     // cmd_xbar_demux_010:src12_valid -> cmd_xbar_mux_057:sink1_valid
	wire         cmd_xbar_demux_010_src12_startofpacket;                                                             // cmd_xbar_demux_010:src12_startofpacket -> cmd_xbar_mux_057:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src12_data;                                                                      // cmd_xbar_demux_010:src12_data -> cmd_xbar_mux_057:sink1_data
	wire  [65:0] cmd_xbar_demux_010_src12_channel;                                                                   // cmd_xbar_demux_010:src12_channel -> cmd_xbar_mux_057:sink1_channel
	wire         cmd_xbar_demux_010_src12_ready;                                                                     // cmd_xbar_mux_057:sink1_ready -> cmd_xbar_demux_010:src12_ready
	wire         cmd_xbar_demux_010_src13_endofpacket;                                                               // cmd_xbar_demux_010:src13_endofpacket -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_010_src13_valid;                                                                     // cmd_xbar_demux_010:src13_valid -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_010_src13_startofpacket;                                                             // cmd_xbar_demux_010:src13_startofpacket -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src13_data;                                                                      // cmd_xbar_demux_010:src13_data -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_010_src13_channel;                                                                   // cmd_xbar_demux_010:src13_channel -> data_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_010_src14_endofpacket;                                                               // cmd_xbar_demux_010:src14_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_010_src14_valid;                                                                     // cmd_xbar_demux_010:src14_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_010_src14_startofpacket;                                                             // cmd_xbar_demux_010:src14_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src14_data;                                                                      // cmd_xbar_demux_010:src14_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_010_src14_channel;                                                                   // cmd_xbar_demux_010:src14_channel -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_010_src15_endofpacket;                                                               // cmd_xbar_demux_010:src15_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_010_src15_valid;                                                                     // cmd_xbar_demux_010:src15_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_010_src15_startofpacket;                                                             // cmd_xbar_demux_010:src15_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src15_data;                                                                      // cmd_xbar_demux_010:src15_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_010_src15_channel;                                                                   // cmd_xbar_demux_010:src15_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_010_src16_endofpacket;                                                               // cmd_xbar_demux_010:src16_endofpacket -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_010_src16_valid;                                                                     // cmd_xbar_demux_010:src16_valid -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_010_src16_startofpacket;                                                             // cmd_xbar_demux_010:src16_startofpacket -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_010_src16_data;                                                                      // cmd_xbar_demux_010:src16_data -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_010_src16_channel;                                                                   // cmd_xbar_demux_010:src16_channel -> high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_011_src0_endofpacket;                                                                // cmd_xbar_demux_011:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_011_src0_valid;                                                                      // cmd_xbar_demux_011:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_011_src0_startofpacket;                                                              // cmd_xbar_demux_011:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src0_data;                                                                       // cmd_xbar_demux_011:src0_data -> cmd_xbar_mux:sink1_data
	wire  [65:0] cmd_xbar_demux_011_src0_channel;                                                                    // cmd_xbar_demux_011:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_011_src0_ready;                                                                      // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_011:src0_ready
	wire         cmd_xbar_demux_011_src1_endofpacket;                                                                // cmd_xbar_demux_011:src1_endofpacket -> cmd_xbar_mux_002:sink3_endofpacket
	wire         cmd_xbar_demux_011_src1_valid;                                                                      // cmd_xbar_demux_011:src1_valid -> cmd_xbar_mux_002:sink3_valid
	wire         cmd_xbar_demux_011_src1_startofpacket;                                                              // cmd_xbar_demux_011:src1_startofpacket -> cmd_xbar_mux_002:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src1_data;                                                                       // cmd_xbar_demux_011:src1_data -> cmd_xbar_mux_002:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src1_channel;                                                                    // cmd_xbar_demux_011:src1_channel -> cmd_xbar_mux_002:sink3_channel
	wire         cmd_xbar_demux_011_src1_ready;                                                                      // cmd_xbar_mux_002:sink3_ready -> cmd_xbar_demux_011:src1_ready
	wire         cmd_xbar_demux_011_src2_endofpacket;                                                                // cmd_xbar_demux_011:src2_endofpacket -> cmd_xbar_mux_003:sink3_endofpacket
	wire         cmd_xbar_demux_011_src2_valid;                                                                      // cmd_xbar_demux_011:src2_valid -> cmd_xbar_mux_003:sink3_valid
	wire         cmd_xbar_demux_011_src2_startofpacket;                                                              // cmd_xbar_demux_011:src2_startofpacket -> cmd_xbar_mux_003:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src2_data;                                                                       // cmd_xbar_demux_011:src2_data -> cmd_xbar_mux_003:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src2_channel;                                                                    // cmd_xbar_demux_011:src2_channel -> cmd_xbar_mux_003:sink3_channel
	wire         cmd_xbar_demux_011_src2_ready;                                                                      // cmd_xbar_mux_003:sink3_ready -> cmd_xbar_demux_011:src2_ready
	wire         cmd_xbar_demux_011_src3_endofpacket;                                                                // cmd_xbar_demux_011:src3_endofpacket -> cmd_xbar_mux_004:sink3_endofpacket
	wire         cmd_xbar_demux_011_src3_valid;                                                                      // cmd_xbar_demux_011:src3_valid -> cmd_xbar_mux_004:sink3_valid
	wire         cmd_xbar_demux_011_src3_startofpacket;                                                              // cmd_xbar_demux_011:src3_startofpacket -> cmd_xbar_mux_004:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src3_data;                                                                       // cmd_xbar_demux_011:src3_data -> cmd_xbar_mux_004:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src3_channel;                                                                    // cmd_xbar_demux_011:src3_channel -> cmd_xbar_mux_004:sink3_channel
	wire         cmd_xbar_demux_011_src3_ready;                                                                      // cmd_xbar_mux_004:sink3_ready -> cmd_xbar_demux_011:src3_ready
	wire         cmd_xbar_demux_011_src4_endofpacket;                                                                // cmd_xbar_demux_011:src4_endofpacket -> cmd_xbar_mux_005:sink3_endofpacket
	wire         cmd_xbar_demux_011_src4_valid;                                                                      // cmd_xbar_demux_011:src4_valid -> cmd_xbar_mux_005:sink3_valid
	wire         cmd_xbar_demux_011_src4_startofpacket;                                                              // cmd_xbar_demux_011:src4_startofpacket -> cmd_xbar_mux_005:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src4_data;                                                                       // cmd_xbar_demux_011:src4_data -> cmd_xbar_mux_005:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src4_channel;                                                                    // cmd_xbar_demux_011:src4_channel -> cmd_xbar_mux_005:sink3_channel
	wire         cmd_xbar_demux_011_src4_ready;                                                                      // cmd_xbar_mux_005:sink3_ready -> cmd_xbar_demux_011:src4_ready
	wire         cmd_xbar_demux_011_src5_endofpacket;                                                                // cmd_xbar_demux_011:src5_endofpacket -> cmd_xbar_mux_006:sink3_endofpacket
	wire         cmd_xbar_demux_011_src5_valid;                                                                      // cmd_xbar_demux_011:src5_valid -> cmd_xbar_mux_006:sink3_valid
	wire         cmd_xbar_demux_011_src5_startofpacket;                                                              // cmd_xbar_demux_011:src5_startofpacket -> cmd_xbar_mux_006:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src5_data;                                                                       // cmd_xbar_demux_011:src5_data -> cmd_xbar_mux_006:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src5_channel;                                                                    // cmd_xbar_demux_011:src5_channel -> cmd_xbar_mux_006:sink3_channel
	wire         cmd_xbar_demux_011_src5_ready;                                                                      // cmd_xbar_mux_006:sink3_ready -> cmd_xbar_demux_011:src5_ready
	wire         cmd_xbar_demux_011_src6_endofpacket;                                                                // cmd_xbar_demux_011:src6_endofpacket -> cmd_xbar_mux_007:sink3_endofpacket
	wire         cmd_xbar_demux_011_src6_valid;                                                                      // cmd_xbar_demux_011:src6_valid -> cmd_xbar_mux_007:sink3_valid
	wire         cmd_xbar_demux_011_src6_startofpacket;                                                              // cmd_xbar_demux_011:src6_startofpacket -> cmd_xbar_mux_007:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src6_data;                                                                       // cmd_xbar_demux_011:src6_data -> cmd_xbar_mux_007:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src6_channel;                                                                    // cmd_xbar_demux_011:src6_channel -> cmd_xbar_mux_007:sink3_channel
	wire         cmd_xbar_demux_011_src6_ready;                                                                      // cmd_xbar_mux_007:sink3_ready -> cmd_xbar_demux_011:src6_ready
	wire         cmd_xbar_demux_011_src7_endofpacket;                                                                // cmd_xbar_demux_011:src7_endofpacket -> cmd_xbar_mux_008:sink3_endofpacket
	wire         cmd_xbar_demux_011_src7_valid;                                                                      // cmd_xbar_demux_011:src7_valid -> cmd_xbar_mux_008:sink3_valid
	wire         cmd_xbar_demux_011_src7_startofpacket;                                                              // cmd_xbar_demux_011:src7_startofpacket -> cmd_xbar_mux_008:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src7_data;                                                                       // cmd_xbar_demux_011:src7_data -> cmd_xbar_mux_008:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src7_channel;                                                                    // cmd_xbar_demux_011:src7_channel -> cmd_xbar_mux_008:sink3_channel
	wire         cmd_xbar_demux_011_src7_ready;                                                                      // cmd_xbar_mux_008:sink3_ready -> cmd_xbar_demux_011:src7_ready
	wire         cmd_xbar_demux_011_src8_endofpacket;                                                                // cmd_xbar_demux_011:src8_endofpacket -> cmd_xbar_mux_009:sink3_endofpacket
	wire         cmd_xbar_demux_011_src8_valid;                                                                      // cmd_xbar_demux_011:src8_valid -> cmd_xbar_mux_009:sink3_valid
	wire         cmd_xbar_demux_011_src8_startofpacket;                                                              // cmd_xbar_demux_011:src8_startofpacket -> cmd_xbar_mux_009:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src8_data;                                                                       // cmd_xbar_demux_011:src8_data -> cmd_xbar_mux_009:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src8_channel;                                                                    // cmd_xbar_demux_011:src8_channel -> cmd_xbar_mux_009:sink3_channel
	wire         cmd_xbar_demux_011_src8_ready;                                                                      // cmd_xbar_mux_009:sink3_ready -> cmd_xbar_demux_011:src8_ready
	wire         cmd_xbar_demux_011_src9_endofpacket;                                                                // cmd_xbar_demux_011:src9_endofpacket -> cmd_xbar_mux_010:sink3_endofpacket
	wire         cmd_xbar_demux_011_src9_valid;                                                                      // cmd_xbar_demux_011:src9_valid -> cmd_xbar_mux_010:sink3_valid
	wire         cmd_xbar_demux_011_src9_startofpacket;                                                              // cmd_xbar_demux_011:src9_startofpacket -> cmd_xbar_mux_010:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src9_data;                                                                       // cmd_xbar_demux_011:src9_data -> cmd_xbar_mux_010:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src9_channel;                                                                    // cmd_xbar_demux_011:src9_channel -> cmd_xbar_mux_010:sink3_channel
	wire         cmd_xbar_demux_011_src9_ready;                                                                      // cmd_xbar_mux_010:sink3_ready -> cmd_xbar_demux_011:src9_ready
	wire         cmd_xbar_demux_011_src10_endofpacket;                                                               // cmd_xbar_demux_011:src10_endofpacket -> cmd_xbar_mux_011:sink3_endofpacket
	wire         cmd_xbar_demux_011_src10_valid;                                                                     // cmd_xbar_demux_011:src10_valid -> cmd_xbar_mux_011:sink3_valid
	wire         cmd_xbar_demux_011_src10_startofpacket;                                                             // cmd_xbar_demux_011:src10_startofpacket -> cmd_xbar_mux_011:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src10_data;                                                                      // cmd_xbar_demux_011:src10_data -> cmd_xbar_mux_011:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src10_channel;                                                                   // cmd_xbar_demux_011:src10_channel -> cmd_xbar_mux_011:sink3_channel
	wire         cmd_xbar_demux_011_src10_ready;                                                                     // cmd_xbar_mux_011:sink3_ready -> cmd_xbar_demux_011:src10_ready
	wire         cmd_xbar_demux_011_src11_endofpacket;                                                               // cmd_xbar_demux_011:src11_endofpacket -> cmd_xbar_mux_012:sink3_endofpacket
	wire         cmd_xbar_demux_011_src11_valid;                                                                     // cmd_xbar_demux_011:src11_valid -> cmd_xbar_mux_012:sink3_valid
	wire         cmd_xbar_demux_011_src11_startofpacket;                                                             // cmd_xbar_demux_011:src11_startofpacket -> cmd_xbar_mux_012:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src11_data;                                                                      // cmd_xbar_demux_011:src11_data -> cmd_xbar_mux_012:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src11_channel;                                                                   // cmd_xbar_demux_011:src11_channel -> cmd_xbar_mux_012:sink3_channel
	wire         cmd_xbar_demux_011_src11_ready;                                                                     // cmd_xbar_mux_012:sink3_ready -> cmd_xbar_demux_011:src11_ready
	wire         cmd_xbar_demux_011_src12_endofpacket;                                                               // cmd_xbar_demux_011:src12_endofpacket -> cmd_xbar_mux_013:sink3_endofpacket
	wire         cmd_xbar_demux_011_src12_valid;                                                                     // cmd_xbar_demux_011:src12_valid -> cmd_xbar_mux_013:sink3_valid
	wire         cmd_xbar_demux_011_src12_startofpacket;                                                             // cmd_xbar_demux_011:src12_startofpacket -> cmd_xbar_mux_013:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src12_data;                                                                      // cmd_xbar_demux_011:src12_data -> cmd_xbar_mux_013:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src12_channel;                                                                   // cmd_xbar_demux_011:src12_channel -> cmd_xbar_mux_013:sink3_channel
	wire         cmd_xbar_demux_011_src12_ready;                                                                     // cmd_xbar_mux_013:sink3_ready -> cmd_xbar_demux_011:src12_ready
	wire         cmd_xbar_demux_011_src13_endofpacket;                                                               // cmd_xbar_demux_011:src13_endofpacket -> cmd_xbar_mux_014:sink3_endofpacket
	wire         cmd_xbar_demux_011_src13_valid;                                                                     // cmd_xbar_demux_011:src13_valid -> cmd_xbar_mux_014:sink3_valid
	wire         cmd_xbar_demux_011_src13_startofpacket;                                                             // cmd_xbar_demux_011:src13_startofpacket -> cmd_xbar_mux_014:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src13_data;                                                                      // cmd_xbar_demux_011:src13_data -> cmd_xbar_mux_014:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src13_channel;                                                                   // cmd_xbar_demux_011:src13_channel -> cmd_xbar_mux_014:sink3_channel
	wire         cmd_xbar_demux_011_src13_ready;                                                                     // cmd_xbar_mux_014:sink3_ready -> cmd_xbar_demux_011:src13_ready
	wire         cmd_xbar_demux_011_src14_endofpacket;                                                               // cmd_xbar_demux_011:src14_endofpacket -> cmd_xbar_mux_015:sink3_endofpacket
	wire         cmd_xbar_demux_011_src14_valid;                                                                     // cmd_xbar_demux_011:src14_valid -> cmd_xbar_mux_015:sink3_valid
	wire         cmd_xbar_demux_011_src14_startofpacket;                                                             // cmd_xbar_demux_011:src14_startofpacket -> cmd_xbar_mux_015:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src14_data;                                                                      // cmd_xbar_demux_011:src14_data -> cmd_xbar_mux_015:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src14_channel;                                                                   // cmd_xbar_demux_011:src14_channel -> cmd_xbar_mux_015:sink3_channel
	wire         cmd_xbar_demux_011_src14_ready;                                                                     // cmd_xbar_mux_015:sink3_ready -> cmd_xbar_demux_011:src14_ready
	wire         cmd_xbar_demux_011_src15_endofpacket;                                                               // cmd_xbar_demux_011:src15_endofpacket -> cmd_xbar_mux_016:sink3_endofpacket
	wire         cmd_xbar_demux_011_src15_valid;                                                                     // cmd_xbar_demux_011:src15_valid -> cmd_xbar_mux_016:sink3_valid
	wire         cmd_xbar_demux_011_src15_startofpacket;                                                             // cmd_xbar_demux_011:src15_startofpacket -> cmd_xbar_mux_016:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src15_data;                                                                      // cmd_xbar_demux_011:src15_data -> cmd_xbar_mux_016:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src15_channel;                                                                   // cmd_xbar_demux_011:src15_channel -> cmd_xbar_mux_016:sink3_channel
	wire         cmd_xbar_demux_011_src15_ready;                                                                     // cmd_xbar_mux_016:sink3_ready -> cmd_xbar_demux_011:src15_ready
	wire         cmd_xbar_demux_011_src16_endofpacket;                                                               // cmd_xbar_demux_011:src16_endofpacket -> cmd_xbar_mux_017:sink3_endofpacket
	wire         cmd_xbar_demux_011_src16_valid;                                                                     // cmd_xbar_demux_011:src16_valid -> cmd_xbar_mux_017:sink3_valid
	wire         cmd_xbar_demux_011_src16_startofpacket;                                                             // cmd_xbar_demux_011:src16_startofpacket -> cmd_xbar_mux_017:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src16_data;                                                                      // cmd_xbar_demux_011:src16_data -> cmd_xbar_mux_017:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src16_channel;                                                                   // cmd_xbar_demux_011:src16_channel -> cmd_xbar_mux_017:sink3_channel
	wire         cmd_xbar_demux_011_src16_ready;                                                                     // cmd_xbar_mux_017:sink3_ready -> cmd_xbar_demux_011:src16_ready
	wire         cmd_xbar_demux_011_src17_endofpacket;                                                               // cmd_xbar_demux_011:src17_endofpacket -> cmd_xbar_mux_018:sink3_endofpacket
	wire         cmd_xbar_demux_011_src17_valid;                                                                     // cmd_xbar_demux_011:src17_valid -> cmd_xbar_mux_018:sink3_valid
	wire         cmd_xbar_demux_011_src17_startofpacket;                                                             // cmd_xbar_demux_011:src17_startofpacket -> cmd_xbar_mux_018:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src17_data;                                                                      // cmd_xbar_demux_011:src17_data -> cmd_xbar_mux_018:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src17_channel;                                                                   // cmd_xbar_demux_011:src17_channel -> cmd_xbar_mux_018:sink3_channel
	wire         cmd_xbar_demux_011_src17_ready;                                                                     // cmd_xbar_mux_018:sink3_ready -> cmd_xbar_demux_011:src17_ready
	wire         cmd_xbar_demux_011_src18_endofpacket;                                                               // cmd_xbar_demux_011:src18_endofpacket -> cmd_xbar_mux_019:sink3_endofpacket
	wire         cmd_xbar_demux_011_src18_valid;                                                                     // cmd_xbar_demux_011:src18_valid -> cmd_xbar_mux_019:sink3_valid
	wire         cmd_xbar_demux_011_src18_startofpacket;                                                             // cmd_xbar_demux_011:src18_startofpacket -> cmd_xbar_mux_019:sink3_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src18_data;                                                                      // cmd_xbar_demux_011:src18_data -> cmd_xbar_mux_019:sink3_data
	wire  [65:0] cmd_xbar_demux_011_src18_channel;                                                                   // cmd_xbar_demux_011:src18_channel -> cmd_xbar_mux_019:sink3_channel
	wire         cmd_xbar_demux_011_src18_ready;                                                                     // cmd_xbar_mux_019:sink3_ready -> cmd_xbar_demux_011:src18_ready
	wire         cmd_xbar_demux_011_src19_endofpacket;                                                               // cmd_xbar_demux_011:src19_endofpacket -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_011_src19_valid;                                                                     // cmd_xbar_demux_011:src19_valid -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_011_src19_startofpacket;                                                             // cmd_xbar_demux_011:src19_startofpacket -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src19_data;                                                                      // cmd_xbar_demux_011:src19_data -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_011_src19_channel;                                                                   // cmd_xbar_demux_011:src19_channel -> data_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_011_src20_endofpacket;                                                               // cmd_xbar_demux_011:src20_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_011_src20_valid;                                                                     // cmd_xbar_demux_011:src20_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_011_src20_startofpacket;                                                             // cmd_xbar_demux_011:src20_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src20_data;                                                                      // cmd_xbar_demux_011:src20_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_011_src20_channel;                                                                   // cmd_xbar_demux_011:src20_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_011_src21_endofpacket;                                                               // cmd_xbar_demux_011:src21_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_011_src21_valid;                                                                     // cmd_xbar_demux_011:src21_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_011_src21_startofpacket;                                                             // cmd_xbar_demux_011:src21_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src21_data;                                                                      // cmd_xbar_demux_011:src21_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_011_src21_channel;                                                                   // cmd_xbar_demux_011:src21_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_011_src22_endofpacket;                                                               // cmd_xbar_demux_011:src22_endofpacket -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_011_src22_valid;                                                                     // cmd_xbar_demux_011:src22_valid -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_011_src22_startofpacket;                                                             // cmd_xbar_demux_011:src22_startofpacket -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_demux_011_src22_data;                                                                      // cmd_xbar_demux_011:src22_data -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_demux_011_src22_channel;                                                                   // cmd_xbar_demux_011:src22_channel -> high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                    // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                          // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                  // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_src0_data;                                                                           // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [65:0] rsp_xbar_demux_src0_channel;                                                                        // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                          // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                    // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_011:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                          // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_011:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                  // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_011:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_src1_data;                                                                           // rsp_xbar_demux:src1_data -> rsp_xbar_mux_011:sink0_data
	wire  [65:0] rsp_xbar_demux_src1_channel;                                                                        // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_011:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                          // rsp_xbar_mux_011:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                      // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                              // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_001_src0_data;                                                                       // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [65:0] rsp_xbar_demux_001_src0_channel;                                                                    // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                      // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                      // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                              // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_002_src0_data;                                                                       // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [65:0] rsp_xbar_demux_002_src0_channel;                                                                    // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                      // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_009:sink0_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                      // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_009:sink0_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                              // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_009:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_002_src1_data;                                                                       // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_009:sink0_data
	wire  [65:0] rsp_xbar_demux_002_src1_channel;                                                                    // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_009:sink0_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                      // rsp_xbar_mux_009:sink0_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_002_src2_endofpacket;                                                                // rsp_xbar_demux_002:src2_endofpacket -> rsp_xbar_mux_010:sink0_endofpacket
	wire         rsp_xbar_demux_002_src2_valid;                                                                      // rsp_xbar_demux_002:src2_valid -> rsp_xbar_mux_010:sink0_valid
	wire         rsp_xbar_demux_002_src2_startofpacket;                                                              // rsp_xbar_demux_002:src2_startofpacket -> rsp_xbar_mux_010:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_002_src2_data;                                                                       // rsp_xbar_demux_002:src2_data -> rsp_xbar_mux_010:sink0_data
	wire  [65:0] rsp_xbar_demux_002_src2_channel;                                                                    // rsp_xbar_demux_002:src2_channel -> rsp_xbar_mux_010:sink0_channel
	wire         rsp_xbar_demux_002_src2_ready;                                                                      // rsp_xbar_mux_010:sink0_ready -> rsp_xbar_demux_002:src2_ready
	wire         rsp_xbar_demux_002_src3_endofpacket;                                                                // rsp_xbar_demux_002:src3_endofpacket -> rsp_xbar_mux_011:sink1_endofpacket
	wire         rsp_xbar_demux_002_src3_valid;                                                                      // rsp_xbar_demux_002:src3_valid -> rsp_xbar_mux_011:sink1_valid
	wire         rsp_xbar_demux_002_src3_startofpacket;                                                              // rsp_xbar_demux_002:src3_startofpacket -> rsp_xbar_mux_011:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_002_src3_data;                                                                       // rsp_xbar_demux_002:src3_data -> rsp_xbar_mux_011:sink1_data
	wire  [65:0] rsp_xbar_demux_002_src3_channel;                                                                    // rsp_xbar_demux_002:src3_channel -> rsp_xbar_mux_011:sink1_channel
	wire         rsp_xbar_demux_002_src3_ready;                                                                      // rsp_xbar_mux_011:sink1_ready -> rsp_xbar_demux_002:src3_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                      // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                              // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_003_src0_data;                                                                       // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire  [65:0] rsp_xbar_demux_003_src0_channel;                                                                    // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                      // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                                // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_009:sink1_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                      // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_009:sink1_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                              // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_009:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_003_src1_data;                                                                       // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_009:sink1_data
	wire  [65:0] rsp_xbar_demux_003_src1_channel;                                                                    // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_009:sink1_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                      // rsp_xbar_mux_009:sink1_ready -> rsp_xbar_demux_003:src1_ready
	wire         rsp_xbar_demux_003_src2_endofpacket;                                                                // rsp_xbar_demux_003:src2_endofpacket -> rsp_xbar_mux_010:sink1_endofpacket
	wire         rsp_xbar_demux_003_src2_valid;                                                                      // rsp_xbar_demux_003:src2_valid -> rsp_xbar_mux_010:sink1_valid
	wire         rsp_xbar_demux_003_src2_startofpacket;                                                              // rsp_xbar_demux_003:src2_startofpacket -> rsp_xbar_mux_010:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_003_src2_data;                                                                       // rsp_xbar_demux_003:src2_data -> rsp_xbar_mux_010:sink1_data
	wire  [65:0] rsp_xbar_demux_003_src2_channel;                                                                    // rsp_xbar_demux_003:src2_channel -> rsp_xbar_mux_010:sink1_channel
	wire         rsp_xbar_demux_003_src2_ready;                                                                      // rsp_xbar_mux_010:sink1_ready -> rsp_xbar_demux_003:src2_ready
	wire         rsp_xbar_demux_003_src3_endofpacket;                                                                // rsp_xbar_demux_003:src3_endofpacket -> rsp_xbar_mux_011:sink2_endofpacket
	wire         rsp_xbar_demux_003_src3_valid;                                                                      // rsp_xbar_demux_003:src3_valid -> rsp_xbar_mux_011:sink2_valid
	wire         rsp_xbar_demux_003_src3_startofpacket;                                                              // rsp_xbar_demux_003:src3_startofpacket -> rsp_xbar_mux_011:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_003_src3_data;                                                                       // rsp_xbar_demux_003:src3_data -> rsp_xbar_mux_011:sink2_data
	wire  [65:0] rsp_xbar_demux_003_src3_channel;                                                                    // rsp_xbar_demux_003:src3_channel -> rsp_xbar_mux_011:sink2_channel
	wire         rsp_xbar_demux_003_src3_ready;                                                                      // rsp_xbar_mux_011:sink2_ready -> rsp_xbar_demux_003:src3_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                      // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                              // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_004_src0_data;                                                                       // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire  [65:0] rsp_xbar_demux_004_src0_channel;                                                                    // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                      // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_004_src1_endofpacket;                                                                // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_009:sink2_endofpacket
	wire         rsp_xbar_demux_004_src1_valid;                                                                      // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_009:sink2_valid
	wire         rsp_xbar_demux_004_src1_startofpacket;                                                              // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_009:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_004_src1_data;                                                                       // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_009:sink2_data
	wire  [65:0] rsp_xbar_demux_004_src1_channel;                                                                    // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_009:sink2_channel
	wire         rsp_xbar_demux_004_src1_ready;                                                                      // rsp_xbar_mux_009:sink2_ready -> rsp_xbar_demux_004:src1_ready
	wire         rsp_xbar_demux_004_src2_endofpacket;                                                                // rsp_xbar_demux_004:src2_endofpacket -> rsp_xbar_mux_010:sink2_endofpacket
	wire         rsp_xbar_demux_004_src2_valid;                                                                      // rsp_xbar_demux_004:src2_valid -> rsp_xbar_mux_010:sink2_valid
	wire         rsp_xbar_demux_004_src2_startofpacket;                                                              // rsp_xbar_demux_004:src2_startofpacket -> rsp_xbar_mux_010:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_004_src2_data;                                                                       // rsp_xbar_demux_004:src2_data -> rsp_xbar_mux_010:sink2_data
	wire  [65:0] rsp_xbar_demux_004_src2_channel;                                                                    // rsp_xbar_demux_004:src2_channel -> rsp_xbar_mux_010:sink2_channel
	wire         rsp_xbar_demux_004_src2_ready;                                                                      // rsp_xbar_mux_010:sink2_ready -> rsp_xbar_demux_004:src2_ready
	wire         rsp_xbar_demux_004_src3_endofpacket;                                                                // rsp_xbar_demux_004:src3_endofpacket -> rsp_xbar_mux_011:sink3_endofpacket
	wire         rsp_xbar_demux_004_src3_valid;                                                                      // rsp_xbar_demux_004:src3_valid -> rsp_xbar_mux_011:sink3_valid
	wire         rsp_xbar_demux_004_src3_startofpacket;                                                              // rsp_xbar_demux_004:src3_startofpacket -> rsp_xbar_mux_011:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_004_src3_data;                                                                       // rsp_xbar_demux_004:src3_data -> rsp_xbar_mux_011:sink3_data
	wire  [65:0] rsp_xbar_demux_004_src3_channel;                                                                    // rsp_xbar_demux_004:src3_channel -> rsp_xbar_mux_011:sink3_channel
	wire         rsp_xbar_demux_004_src3_ready;                                                                      // rsp_xbar_mux_011:sink3_ready -> rsp_xbar_demux_004:src3_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                      // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                              // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_005_src0_data;                                                                       // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire  [65:0] rsp_xbar_demux_005_src0_channel;                                                                    // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                      // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_005_src1_endofpacket;                                                                // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_009:sink3_endofpacket
	wire         rsp_xbar_demux_005_src1_valid;                                                                      // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_009:sink3_valid
	wire         rsp_xbar_demux_005_src1_startofpacket;                                                              // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_009:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_005_src1_data;                                                                       // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_009:sink3_data
	wire  [65:0] rsp_xbar_demux_005_src1_channel;                                                                    // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_009:sink3_channel
	wire         rsp_xbar_demux_005_src1_ready;                                                                      // rsp_xbar_mux_009:sink3_ready -> rsp_xbar_demux_005:src1_ready
	wire         rsp_xbar_demux_005_src2_endofpacket;                                                                // rsp_xbar_demux_005:src2_endofpacket -> rsp_xbar_mux_010:sink3_endofpacket
	wire         rsp_xbar_demux_005_src2_valid;                                                                      // rsp_xbar_demux_005:src2_valid -> rsp_xbar_mux_010:sink3_valid
	wire         rsp_xbar_demux_005_src2_startofpacket;                                                              // rsp_xbar_demux_005:src2_startofpacket -> rsp_xbar_mux_010:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_005_src2_data;                                                                       // rsp_xbar_demux_005:src2_data -> rsp_xbar_mux_010:sink3_data
	wire  [65:0] rsp_xbar_demux_005_src2_channel;                                                                    // rsp_xbar_demux_005:src2_channel -> rsp_xbar_mux_010:sink3_channel
	wire         rsp_xbar_demux_005_src2_ready;                                                                      // rsp_xbar_mux_010:sink3_ready -> rsp_xbar_demux_005:src2_ready
	wire         rsp_xbar_demux_005_src3_endofpacket;                                                                // rsp_xbar_demux_005:src3_endofpacket -> rsp_xbar_mux_011:sink4_endofpacket
	wire         rsp_xbar_demux_005_src3_valid;                                                                      // rsp_xbar_demux_005:src3_valid -> rsp_xbar_mux_011:sink4_valid
	wire         rsp_xbar_demux_005_src3_startofpacket;                                                              // rsp_xbar_demux_005:src3_startofpacket -> rsp_xbar_mux_011:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_005_src3_data;                                                                       // rsp_xbar_demux_005:src3_data -> rsp_xbar_mux_011:sink4_data
	wire  [65:0] rsp_xbar_demux_005_src3_channel;                                                                    // rsp_xbar_demux_005:src3_channel -> rsp_xbar_mux_011:sink4_channel
	wire         rsp_xbar_demux_005_src3_ready;                                                                      // rsp_xbar_mux_011:sink4_ready -> rsp_xbar_demux_005:src3_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                      // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                              // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_006_src0_data;                                                                       // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire  [65:0] rsp_xbar_demux_006_src0_channel;                                                                    // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                      // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_006_src1_endofpacket;                                                                // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_009:sink4_endofpacket
	wire         rsp_xbar_demux_006_src1_valid;                                                                      // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_009:sink4_valid
	wire         rsp_xbar_demux_006_src1_startofpacket;                                                              // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_009:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_006_src1_data;                                                                       // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_009:sink4_data
	wire  [65:0] rsp_xbar_demux_006_src1_channel;                                                                    // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_009:sink4_channel
	wire         rsp_xbar_demux_006_src1_ready;                                                                      // rsp_xbar_mux_009:sink4_ready -> rsp_xbar_demux_006:src1_ready
	wire         rsp_xbar_demux_006_src2_endofpacket;                                                                // rsp_xbar_demux_006:src2_endofpacket -> rsp_xbar_mux_010:sink4_endofpacket
	wire         rsp_xbar_demux_006_src2_valid;                                                                      // rsp_xbar_demux_006:src2_valid -> rsp_xbar_mux_010:sink4_valid
	wire         rsp_xbar_demux_006_src2_startofpacket;                                                              // rsp_xbar_demux_006:src2_startofpacket -> rsp_xbar_mux_010:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_006_src2_data;                                                                       // rsp_xbar_demux_006:src2_data -> rsp_xbar_mux_010:sink4_data
	wire  [65:0] rsp_xbar_demux_006_src2_channel;                                                                    // rsp_xbar_demux_006:src2_channel -> rsp_xbar_mux_010:sink4_channel
	wire         rsp_xbar_demux_006_src2_ready;                                                                      // rsp_xbar_mux_010:sink4_ready -> rsp_xbar_demux_006:src2_ready
	wire         rsp_xbar_demux_006_src3_endofpacket;                                                                // rsp_xbar_demux_006:src3_endofpacket -> rsp_xbar_mux_011:sink5_endofpacket
	wire         rsp_xbar_demux_006_src3_valid;                                                                      // rsp_xbar_demux_006:src3_valid -> rsp_xbar_mux_011:sink5_valid
	wire         rsp_xbar_demux_006_src3_startofpacket;                                                              // rsp_xbar_demux_006:src3_startofpacket -> rsp_xbar_mux_011:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_006_src3_data;                                                                       // rsp_xbar_demux_006:src3_data -> rsp_xbar_mux_011:sink5_data
	wire  [65:0] rsp_xbar_demux_006_src3_channel;                                                                    // rsp_xbar_demux_006:src3_channel -> rsp_xbar_mux_011:sink5_channel
	wire         rsp_xbar_demux_006_src3_ready;                                                                      // rsp_xbar_mux_011:sink5_ready -> rsp_xbar_demux_006:src3_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                      // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                              // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_007_src0_data;                                                                       // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire  [65:0] rsp_xbar_demux_007_src0_channel;                                                                    // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                      // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_007_src1_endofpacket;                                                                // rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_009:sink5_endofpacket
	wire         rsp_xbar_demux_007_src1_valid;                                                                      // rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_009:sink5_valid
	wire         rsp_xbar_demux_007_src1_startofpacket;                                                              // rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_009:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_007_src1_data;                                                                       // rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_009:sink5_data
	wire  [65:0] rsp_xbar_demux_007_src1_channel;                                                                    // rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_009:sink5_channel
	wire         rsp_xbar_demux_007_src1_ready;                                                                      // rsp_xbar_mux_009:sink5_ready -> rsp_xbar_demux_007:src1_ready
	wire         rsp_xbar_demux_007_src2_endofpacket;                                                                // rsp_xbar_demux_007:src2_endofpacket -> rsp_xbar_mux_010:sink5_endofpacket
	wire         rsp_xbar_demux_007_src2_valid;                                                                      // rsp_xbar_demux_007:src2_valid -> rsp_xbar_mux_010:sink5_valid
	wire         rsp_xbar_demux_007_src2_startofpacket;                                                              // rsp_xbar_demux_007:src2_startofpacket -> rsp_xbar_mux_010:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_007_src2_data;                                                                       // rsp_xbar_demux_007:src2_data -> rsp_xbar_mux_010:sink5_data
	wire  [65:0] rsp_xbar_demux_007_src2_channel;                                                                    // rsp_xbar_demux_007:src2_channel -> rsp_xbar_mux_010:sink5_channel
	wire         rsp_xbar_demux_007_src2_ready;                                                                      // rsp_xbar_mux_010:sink5_ready -> rsp_xbar_demux_007:src2_ready
	wire         rsp_xbar_demux_007_src3_endofpacket;                                                                // rsp_xbar_demux_007:src3_endofpacket -> rsp_xbar_mux_011:sink6_endofpacket
	wire         rsp_xbar_demux_007_src3_valid;                                                                      // rsp_xbar_demux_007:src3_valid -> rsp_xbar_mux_011:sink6_valid
	wire         rsp_xbar_demux_007_src3_startofpacket;                                                              // rsp_xbar_demux_007:src3_startofpacket -> rsp_xbar_mux_011:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_007_src3_data;                                                                       // rsp_xbar_demux_007:src3_data -> rsp_xbar_mux_011:sink6_data
	wire  [65:0] rsp_xbar_demux_007_src3_channel;                                                                    // rsp_xbar_demux_007:src3_channel -> rsp_xbar_mux_011:sink6_channel
	wire         rsp_xbar_demux_007_src3_ready;                                                                      // rsp_xbar_mux_011:sink6_ready -> rsp_xbar_demux_007:src3_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                      // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                              // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_008_src0_data;                                                                       // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire  [65:0] rsp_xbar_demux_008_src0_channel;                                                                    // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                      // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_008_src1_endofpacket;                                                                // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_009:sink6_endofpacket
	wire         rsp_xbar_demux_008_src1_valid;                                                                      // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_009:sink6_valid
	wire         rsp_xbar_demux_008_src1_startofpacket;                                                              // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_009:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_008_src1_data;                                                                       // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_009:sink6_data
	wire  [65:0] rsp_xbar_demux_008_src1_channel;                                                                    // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_009:sink6_channel
	wire         rsp_xbar_demux_008_src1_ready;                                                                      // rsp_xbar_mux_009:sink6_ready -> rsp_xbar_demux_008:src1_ready
	wire         rsp_xbar_demux_008_src2_endofpacket;                                                                // rsp_xbar_demux_008:src2_endofpacket -> rsp_xbar_mux_010:sink6_endofpacket
	wire         rsp_xbar_demux_008_src2_valid;                                                                      // rsp_xbar_demux_008:src2_valid -> rsp_xbar_mux_010:sink6_valid
	wire         rsp_xbar_demux_008_src2_startofpacket;                                                              // rsp_xbar_demux_008:src2_startofpacket -> rsp_xbar_mux_010:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_008_src2_data;                                                                       // rsp_xbar_demux_008:src2_data -> rsp_xbar_mux_010:sink6_data
	wire  [65:0] rsp_xbar_demux_008_src2_channel;                                                                    // rsp_xbar_demux_008:src2_channel -> rsp_xbar_mux_010:sink6_channel
	wire         rsp_xbar_demux_008_src2_ready;                                                                      // rsp_xbar_mux_010:sink6_ready -> rsp_xbar_demux_008:src2_ready
	wire         rsp_xbar_demux_008_src3_endofpacket;                                                                // rsp_xbar_demux_008:src3_endofpacket -> rsp_xbar_mux_011:sink7_endofpacket
	wire         rsp_xbar_demux_008_src3_valid;                                                                      // rsp_xbar_demux_008:src3_valid -> rsp_xbar_mux_011:sink7_valid
	wire         rsp_xbar_demux_008_src3_startofpacket;                                                              // rsp_xbar_demux_008:src3_startofpacket -> rsp_xbar_mux_011:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_008_src3_data;                                                                       // rsp_xbar_demux_008:src3_data -> rsp_xbar_mux_011:sink7_data
	wire  [65:0] rsp_xbar_demux_008_src3_channel;                                                                    // rsp_xbar_demux_008:src3_channel -> rsp_xbar_mux_011:sink7_channel
	wire         rsp_xbar_demux_008_src3_ready;                                                                      // rsp_xbar_mux_011:sink7_ready -> rsp_xbar_demux_008:src3_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                      // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                              // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_009_src0_data;                                                                       // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	wire  [65:0] rsp_xbar_demux_009_src0_channel;                                                                    // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                      // rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_009_src1_endofpacket;                                                                // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_009:sink7_endofpacket
	wire         rsp_xbar_demux_009_src1_valid;                                                                      // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_009:sink7_valid
	wire         rsp_xbar_demux_009_src1_startofpacket;                                                              // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_009:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_009_src1_data;                                                                       // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_009:sink7_data
	wire  [65:0] rsp_xbar_demux_009_src1_channel;                                                                    // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_009:sink7_channel
	wire         rsp_xbar_demux_009_src1_ready;                                                                      // rsp_xbar_mux_009:sink7_ready -> rsp_xbar_demux_009:src1_ready
	wire         rsp_xbar_demux_009_src2_endofpacket;                                                                // rsp_xbar_demux_009:src2_endofpacket -> rsp_xbar_mux_010:sink7_endofpacket
	wire         rsp_xbar_demux_009_src2_valid;                                                                      // rsp_xbar_demux_009:src2_valid -> rsp_xbar_mux_010:sink7_valid
	wire         rsp_xbar_demux_009_src2_startofpacket;                                                              // rsp_xbar_demux_009:src2_startofpacket -> rsp_xbar_mux_010:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_009_src2_data;                                                                       // rsp_xbar_demux_009:src2_data -> rsp_xbar_mux_010:sink7_data
	wire  [65:0] rsp_xbar_demux_009_src2_channel;                                                                    // rsp_xbar_demux_009:src2_channel -> rsp_xbar_mux_010:sink7_channel
	wire         rsp_xbar_demux_009_src2_ready;                                                                      // rsp_xbar_mux_010:sink7_ready -> rsp_xbar_demux_009:src2_ready
	wire         rsp_xbar_demux_009_src3_endofpacket;                                                                // rsp_xbar_demux_009:src3_endofpacket -> rsp_xbar_mux_011:sink8_endofpacket
	wire         rsp_xbar_demux_009_src3_valid;                                                                      // rsp_xbar_demux_009:src3_valid -> rsp_xbar_mux_011:sink8_valid
	wire         rsp_xbar_demux_009_src3_startofpacket;                                                              // rsp_xbar_demux_009:src3_startofpacket -> rsp_xbar_mux_011:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_009_src3_data;                                                                       // rsp_xbar_demux_009:src3_data -> rsp_xbar_mux_011:sink8_data
	wire  [65:0] rsp_xbar_demux_009_src3_channel;                                                                    // rsp_xbar_demux_009:src3_channel -> rsp_xbar_mux_011:sink8_channel
	wire         rsp_xbar_demux_009_src3_ready;                                                                      // rsp_xbar_mux_011:sink8_ready -> rsp_xbar_demux_009:src3_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                      // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                              // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_010_src0_data;                                                                       // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	wire  [65:0] rsp_xbar_demux_010_src0_channel;                                                                    // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                      // rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_010_src1_endofpacket;                                                                // rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_009:sink8_endofpacket
	wire         rsp_xbar_demux_010_src1_valid;                                                                      // rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_009:sink8_valid
	wire         rsp_xbar_demux_010_src1_startofpacket;                                                              // rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_009:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_010_src1_data;                                                                       // rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_009:sink8_data
	wire  [65:0] rsp_xbar_demux_010_src1_channel;                                                                    // rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_009:sink8_channel
	wire         rsp_xbar_demux_010_src1_ready;                                                                      // rsp_xbar_mux_009:sink8_ready -> rsp_xbar_demux_010:src1_ready
	wire         rsp_xbar_demux_010_src2_endofpacket;                                                                // rsp_xbar_demux_010:src2_endofpacket -> rsp_xbar_mux_010:sink8_endofpacket
	wire         rsp_xbar_demux_010_src2_valid;                                                                      // rsp_xbar_demux_010:src2_valid -> rsp_xbar_mux_010:sink8_valid
	wire         rsp_xbar_demux_010_src2_startofpacket;                                                              // rsp_xbar_demux_010:src2_startofpacket -> rsp_xbar_mux_010:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_010_src2_data;                                                                       // rsp_xbar_demux_010:src2_data -> rsp_xbar_mux_010:sink8_data
	wire  [65:0] rsp_xbar_demux_010_src2_channel;                                                                    // rsp_xbar_demux_010:src2_channel -> rsp_xbar_mux_010:sink8_channel
	wire         rsp_xbar_demux_010_src2_ready;                                                                      // rsp_xbar_mux_010:sink8_ready -> rsp_xbar_demux_010:src2_ready
	wire         rsp_xbar_demux_010_src3_endofpacket;                                                                // rsp_xbar_demux_010:src3_endofpacket -> rsp_xbar_mux_011:sink9_endofpacket
	wire         rsp_xbar_demux_010_src3_valid;                                                                      // rsp_xbar_demux_010:src3_valid -> rsp_xbar_mux_011:sink9_valid
	wire         rsp_xbar_demux_010_src3_startofpacket;                                                              // rsp_xbar_demux_010:src3_startofpacket -> rsp_xbar_mux_011:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_010_src3_data;                                                                       // rsp_xbar_demux_010:src3_data -> rsp_xbar_mux_011:sink9_data
	wire  [65:0] rsp_xbar_demux_010_src3_channel;                                                                    // rsp_xbar_demux_010:src3_channel -> rsp_xbar_mux_011:sink9_channel
	wire         rsp_xbar_demux_010_src3_ready;                                                                      // rsp_xbar_mux_011:sink9_ready -> rsp_xbar_demux_010:src3_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                                // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                      // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                              // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	wire  [94:0] rsp_xbar_demux_011_src0_data;                                                                       // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	wire  [65:0] rsp_xbar_demux_011_src0_channel;                                                                    // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                      // rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_011_src1_endofpacket;                                                                // rsp_xbar_demux_011:src1_endofpacket -> rsp_xbar_mux_005:sink0_endofpacket
	wire         rsp_xbar_demux_011_src1_valid;                                                                      // rsp_xbar_demux_011:src1_valid -> rsp_xbar_mux_005:sink0_valid
	wire         rsp_xbar_demux_011_src1_startofpacket;                                                              // rsp_xbar_demux_011:src1_startofpacket -> rsp_xbar_mux_005:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_011_src1_data;                                                                       // rsp_xbar_demux_011:src1_data -> rsp_xbar_mux_005:sink0_data
	wire  [65:0] rsp_xbar_demux_011_src1_channel;                                                                    // rsp_xbar_demux_011:src1_channel -> rsp_xbar_mux_005:sink0_channel
	wire         rsp_xbar_demux_011_src1_ready;                                                                      // rsp_xbar_mux_005:sink0_ready -> rsp_xbar_demux_011:src1_ready
	wire         rsp_xbar_demux_011_src2_endofpacket;                                                                // rsp_xbar_demux_011:src2_endofpacket -> rsp_xbar_mux_006:sink0_endofpacket
	wire         rsp_xbar_demux_011_src2_valid;                                                                      // rsp_xbar_demux_011:src2_valid -> rsp_xbar_mux_006:sink0_valid
	wire         rsp_xbar_demux_011_src2_startofpacket;                                                              // rsp_xbar_demux_011:src2_startofpacket -> rsp_xbar_mux_006:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_011_src2_data;                                                                       // rsp_xbar_demux_011:src2_data -> rsp_xbar_mux_006:sink0_data
	wire  [65:0] rsp_xbar_demux_011_src2_channel;                                                                    // rsp_xbar_demux_011:src2_channel -> rsp_xbar_mux_006:sink0_channel
	wire         rsp_xbar_demux_011_src2_ready;                                                                      // rsp_xbar_mux_006:sink0_ready -> rsp_xbar_demux_011:src2_ready
	wire         rsp_xbar_demux_011_src3_endofpacket;                                                                // rsp_xbar_demux_011:src3_endofpacket -> rsp_xbar_mux_011:sink10_endofpacket
	wire         rsp_xbar_demux_011_src3_valid;                                                                      // rsp_xbar_demux_011:src3_valid -> rsp_xbar_mux_011:sink10_valid
	wire         rsp_xbar_demux_011_src3_startofpacket;                                                              // rsp_xbar_demux_011:src3_startofpacket -> rsp_xbar_mux_011:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_011_src3_data;                                                                       // rsp_xbar_demux_011:src3_data -> rsp_xbar_mux_011:sink10_data
	wire  [65:0] rsp_xbar_demux_011_src3_channel;                                                                    // rsp_xbar_demux_011:src3_channel -> rsp_xbar_mux_011:sink10_channel
	wire         rsp_xbar_demux_011_src3_ready;                                                                      // rsp_xbar_mux_011:sink10_ready -> rsp_xbar_demux_011:src3_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                                // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                      // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                              // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	wire  [94:0] rsp_xbar_demux_012_src0_data;                                                                       // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	wire  [65:0] rsp_xbar_demux_012_src0_channel;                                                                    // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                      // rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_012_src1_endofpacket;                                                                // rsp_xbar_demux_012:src1_endofpacket -> rsp_xbar_mux_005:sink1_endofpacket
	wire         rsp_xbar_demux_012_src1_valid;                                                                      // rsp_xbar_demux_012:src1_valid -> rsp_xbar_mux_005:sink1_valid
	wire         rsp_xbar_demux_012_src1_startofpacket;                                                              // rsp_xbar_demux_012:src1_startofpacket -> rsp_xbar_mux_005:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_012_src1_data;                                                                       // rsp_xbar_demux_012:src1_data -> rsp_xbar_mux_005:sink1_data
	wire  [65:0] rsp_xbar_demux_012_src1_channel;                                                                    // rsp_xbar_demux_012:src1_channel -> rsp_xbar_mux_005:sink1_channel
	wire         rsp_xbar_demux_012_src1_ready;                                                                      // rsp_xbar_mux_005:sink1_ready -> rsp_xbar_demux_012:src1_ready
	wire         rsp_xbar_demux_012_src2_endofpacket;                                                                // rsp_xbar_demux_012:src2_endofpacket -> rsp_xbar_mux_006:sink1_endofpacket
	wire         rsp_xbar_demux_012_src2_valid;                                                                      // rsp_xbar_demux_012:src2_valid -> rsp_xbar_mux_006:sink1_valid
	wire         rsp_xbar_demux_012_src2_startofpacket;                                                              // rsp_xbar_demux_012:src2_startofpacket -> rsp_xbar_mux_006:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_012_src2_data;                                                                       // rsp_xbar_demux_012:src2_data -> rsp_xbar_mux_006:sink1_data
	wire  [65:0] rsp_xbar_demux_012_src2_channel;                                                                    // rsp_xbar_demux_012:src2_channel -> rsp_xbar_mux_006:sink1_channel
	wire         rsp_xbar_demux_012_src2_ready;                                                                      // rsp_xbar_mux_006:sink1_ready -> rsp_xbar_demux_012:src2_ready
	wire         rsp_xbar_demux_012_src3_endofpacket;                                                                // rsp_xbar_demux_012:src3_endofpacket -> rsp_xbar_mux_011:sink11_endofpacket
	wire         rsp_xbar_demux_012_src3_valid;                                                                      // rsp_xbar_demux_012:src3_valid -> rsp_xbar_mux_011:sink11_valid
	wire         rsp_xbar_demux_012_src3_startofpacket;                                                              // rsp_xbar_demux_012:src3_startofpacket -> rsp_xbar_mux_011:sink11_startofpacket
	wire  [94:0] rsp_xbar_demux_012_src3_data;                                                                       // rsp_xbar_demux_012:src3_data -> rsp_xbar_mux_011:sink11_data
	wire  [65:0] rsp_xbar_demux_012_src3_channel;                                                                    // rsp_xbar_demux_012:src3_channel -> rsp_xbar_mux_011:sink11_channel
	wire         rsp_xbar_demux_012_src3_ready;                                                                      // rsp_xbar_mux_011:sink11_ready -> rsp_xbar_demux_012:src3_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                                // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                      // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                              // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	wire  [94:0] rsp_xbar_demux_013_src0_data;                                                                       // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	wire  [65:0] rsp_xbar_demux_013_src0_channel;                                                                    // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                      // rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_013_src1_endofpacket;                                                                // rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_005:sink2_endofpacket
	wire         rsp_xbar_demux_013_src1_valid;                                                                      // rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_005:sink2_valid
	wire         rsp_xbar_demux_013_src1_startofpacket;                                                              // rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_005:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_013_src1_data;                                                                       // rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_005:sink2_data
	wire  [65:0] rsp_xbar_demux_013_src1_channel;                                                                    // rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_005:sink2_channel
	wire         rsp_xbar_demux_013_src1_ready;                                                                      // rsp_xbar_mux_005:sink2_ready -> rsp_xbar_demux_013:src1_ready
	wire         rsp_xbar_demux_013_src2_endofpacket;                                                                // rsp_xbar_demux_013:src2_endofpacket -> rsp_xbar_mux_006:sink2_endofpacket
	wire         rsp_xbar_demux_013_src2_valid;                                                                      // rsp_xbar_demux_013:src2_valid -> rsp_xbar_mux_006:sink2_valid
	wire         rsp_xbar_demux_013_src2_startofpacket;                                                              // rsp_xbar_demux_013:src2_startofpacket -> rsp_xbar_mux_006:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_013_src2_data;                                                                       // rsp_xbar_demux_013:src2_data -> rsp_xbar_mux_006:sink2_data
	wire  [65:0] rsp_xbar_demux_013_src2_channel;                                                                    // rsp_xbar_demux_013:src2_channel -> rsp_xbar_mux_006:sink2_channel
	wire         rsp_xbar_demux_013_src2_ready;                                                                      // rsp_xbar_mux_006:sink2_ready -> rsp_xbar_demux_013:src2_ready
	wire         rsp_xbar_demux_013_src3_endofpacket;                                                                // rsp_xbar_demux_013:src3_endofpacket -> rsp_xbar_mux_011:sink12_endofpacket
	wire         rsp_xbar_demux_013_src3_valid;                                                                      // rsp_xbar_demux_013:src3_valid -> rsp_xbar_mux_011:sink12_valid
	wire         rsp_xbar_demux_013_src3_startofpacket;                                                              // rsp_xbar_demux_013:src3_startofpacket -> rsp_xbar_mux_011:sink12_startofpacket
	wire  [94:0] rsp_xbar_demux_013_src3_data;                                                                       // rsp_xbar_demux_013:src3_data -> rsp_xbar_mux_011:sink12_data
	wire  [65:0] rsp_xbar_demux_013_src3_channel;                                                                    // rsp_xbar_demux_013:src3_channel -> rsp_xbar_mux_011:sink12_channel
	wire         rsp_xbar_demux_013_src3_ready;                                                                      // rsp_xbar_mux_011:sink12_ready -> rsp_xbar_demux_013:src3_ready
	wire         rsp_xbar_demux_014_src0_endofpacket;                                                                // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux:sink14_endofpacket
	wire         rsp_xbar_demux_014_src0_valid;                                                                      // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux:sink14_valid
	wire         rsp_xbar_demux_014_src0_startofpacket;                                                              // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux:sink14_startofpacket
	wire  [94:0] rsp_xbar_demux_014_src0_data;                                                                       // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux:sink14_data
	wire  [65:0] rsp_xbar_demux_014_src0_channel;                                                                    // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux:sink14_channel
	wire         rsp_xbar_demux_014_src0_ready;                                                                      // rsp_xbar_mux:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire         rsp_xbar_demux_014_src1_endofpacket;                                                                // rsp_xbar_demux_014:src1_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire         rsp_xbar_demux_014_src1_valid;                                                                      // rsp_xbar_demux_014:src1_valid -> rsp_xbar_mux_003:sink0_valid
	wire         rsp_xbar_demux_014_src1_startofpacket;                                                              // rsp_xbar_demux_014:src1_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_014_src1_data;                                                                       // rsp_xbar_demux_014:src1_data -> rsp_xbar_mux_003:sink0_data
	wire  [65:0] rsp_xbar_demux_014_src1_channel;                                                                    // rsp_xbar_demux_014:src1_channel -> rsp_xbar_mux_003:sink0_channel
	wire         rsp_xbar_demux_014_src1_ready;                                                                      // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_014:src1_ready
	wire         rsp_xbar_demux_014_src2_endofpacket;                                                                // rsp_xbar_demux_014:src2_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	wire         rsp_xbar_demux_014_src2_valid;                                                                      // rsp_xbar_demux_014:src2_valid -> rsp_xbar_mux_004:sink0_valid
	wire         rsp_xbar_demux_014_src2_startofpacket;                                                              // rsp_xbar_demux_014:src2_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_014_src2_data;                                                                       // rsp_xbar_demux_014:src2_data -> rsp_xbar_mux_004:sink0_data
	wire  [65:0] rsp_xbar_demux_014_src2_channel;                                                                    // rsp_xbar_demux_014:src2_channel -> rsp_xbar_mux_004:sink0_channel
	wire         rsp_xbar_demux_014_src2_ready;                                                                      // rsp_xbar_mux_004:sink0_ready -> rsp_xbar_demux_014:src2_ready
	wire         rsp_xbar_demux_014_src3_endofpacket;                                                                // rsp_xbar_demux_014:src3_endofpacket -> rsp_xbar_mux_011:sink13_endofpacket
	wire         rsp_xbar_demux_014_src3_valid;                                                                      // rsp_xbar_demux_014:src3_valid -> rsp_xbar_mux_011:sink13_valid
	wire         rsp_xbar_demux_014_src3_startofpacket;                                                              // rsp_xbar_demux_014:src3_startofpacket -> rsp_xbar_mux_011:sink13_startofpacket
	wire  [94:0] rsp_xbar_demux_014_src3_data;                                                                       // rsp_xbar_demux_014:src3_data -> rsp_xbar_mux_011:sink13_data
	wire  [65:0] rsp_xbar_demux_014_src3_channel;                                                                    // rsp_xbar_demux_014:src3_channel -> rsp_xbar_mux_011:sink13_channel
	wire         rsp_xbar_demux_014_src3_ready;                                                                      // rsp_xbar_mux_011:sink13_ready -> rsp_xbar_demux_014:src3_ready
	wire         rsp_xbar_demux_015_src0_endofpacket;                                                                // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux:sink15_endofpacket
	wire         rsp_xbar_demux_015_src0_valid;                                                                      // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux:sink15_valid
	wire         rsp_xbar_demux_015_src0_startofpacket;                                                              // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux:sink15_startofpacket
	wire  [94:0] rsp_xbar_demux_015_src0_data;                                                                       // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux:sink15_data
	wire  [65:0] rsp_xbar_demux_015_src0_channel;                                                                    // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux:sink15_channel
	wire         rsp_xbar_demux_015_src0_ready;                                                                      // rsp_xbar_mux:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire         rsp_xbar_demux_015_src1_endofpacket;                                                                // rsp_xbar_demux_015:src1_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire         rsp_xbar_demux_015_src1_valid;                                                                      // rsp_xbar_demux_015:src1_valid -> rsp_xbar_mux_003:sink1_valid
	wire         rsp_xbar_demux_015_src1_startofpacket;                                                              // rsp_xbar_demux_015:src1_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_015_src1_data;                                                                       // rsp_xbar_demux_015:src1_data -> rsp_xbar_mux_003:sink1_data
	wire  [65:0] rsp_xbar_demux_015_src1_channel;                                                                    // rsp_xbar_demux_015:src1_channel -> rsp_xbar_mux_003:sink1_channel
	wire         rsp_xbar_demux_015_src1_ready;                                                                      // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_015:src1_ready
	wire         rsp_xbar_demux_015_src2_endofpacket;                                                                // rsp_xbar_demux_015:src2_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	wire         rsp_xbar_demux_015_src2_valid;                                                                      // rsp_xbar_demux_015:src2_valid -> rsp_xbar_mux_004:sink1_valid
	wire         rsp_xbar_demux_015_src2_startofpacket;                                                              // rsp_xbar_demux_015:src2_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_015_src2_data;                                                                       // rsp_xbar_demux_015:src2_data -> rsp_xbar_mux_004:sink1_data
	wire  [65:0] rsp_xbar_demux_015_src2_channel;                                                                    // rsp_xbar_demux_015:src2_channel -> rsp_xbar_mux_004:sink1_channel
	wire         rsp_xbar_demux_015_src2_ready;                                                                      // rsp_xbar_mux_004:sink1_ready -> rsp_xbar_demux_015:src2_ready
	wire         rsp_xbar_demux_015_src3_endofpacket;                                                                // rsp_xbar_demux_015:src3_endofpacket -> rsp_xbar_mux_011:sink14_endofpacket
	wire         rsp_xbar_demux_015_src3_valid;                                                                      // rsp_xbar_demux_015:src3_valid -> rsp_xbar_mux_011:sink14_valid
	wire         rsp_xbar_demux_015_src3_startofpacket;                                                              // rsp_xbar_demux_015:src3_startofpacket -> rsp_xbar_mux_011:sink14_startofpacket
	wire  [94:0] rsp_xbar_demux_015_src3_data;                                                                       // rsp_xbar_demux_015:src3_data -> rsp_xbar_mux_011:sink14_data
	wire  [65:0] rsp_xbar_demux_015_src3_channel;                                                                    // rsp_xbar_demux_015:src3_channel -> rsp_xbar_mux_011:sink14_channel
	wire         rsp_xbar_demux_015_src3_ready;                                                                      // rsp_xbar_mux_011:sink14_ready -> rsp_xbar_demux_015:src3_ready
	wire         rsp_xbar_demux_016_src0_endofpacket;                                                                // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux:sink16_endofpacket
	wire         rsp_xbar_demux_016_src0_valid;                                                                      // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux:sink16_valid
	wire         rsp_xbar_demux_016_src0_startofpacket;                                                              // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux:sink16_startofpacket
	wire  [94:0] rsp_xbar_demux_016_src0_data;                                                                       // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux:sink16_data
	wire  [65:0] rsp_xbar_demux_016_src0_channel;                                                                    // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux:sink16_channel
	wire         rsp_xbar_demux_016_src0_ready;                                                                      // rsp_xbar_mux:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire         rsp_xbar_demux_016_src1_endofpacket;                                                                // rsp_xbar_demux_016:src1_endofpacket -> rsp_xbar_mux_003:sink2_endofpacket
	wire         rsp_xbar_demux_016_src1_valid;                                                                      // rsp_xbar_demux_016:src1_valid -> rsp_xbar_mux_003:sink2_valid
	wire         rsp_xbar_demux_016_src1_startofpacket;                                                              // rsp_xbar_demux_016:src1_startofpacket -> rsp_xbar_mux_003:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_016_src1_data;                                                                       // rsp_xbar_demux_016:src1_data -> rsp_xbar_mux_003:sink2_data
	wire  [65:0] rsp_xbar_demux_016_src1_channel;                                                                    // rsp_xbar_demux_016:src1_channel -> rsp_xbar_mux_003:sink2_channel
	wire         rsp_xbar_demux_016_src1_ready;                                                                      // rsp_xbar_mux_003:sink2_ready -> rsp_xbar_demux_016:src1_ready
	wire         rsp_xbar_demux_016_src2_endofpacket;                                                                // rsp_xbar_demux_016:src2_endofpacket -> rsp_xbar_mux_004:sink2_endofpacket
	wire         rsp_xbar_demux_016_src2_valid;                                                                      // rsp_xbar_demux_016:src2_valid -> rsp_xbar_mux_004:sink2_valid
	wire         rsp_xbar_demux_016_src2_startofpacket;                                                              // rsp_xbar_demux_016:src2_startofpacket -> rsp_xbar_mux_004:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_016_src2_data;                                                                       // rsp_xbar_demux_016:src2_data -> rsp_xbar_mux_004:sink2_data
	wire  [65:0] rsp_xbar_demux_016_src2_channel;                                                                    // rsp_xbar_demux_016:src2_channel -> rsp_xbar_mux_004:sink2_channel
	wire         rsp_xbar_demux_016_src2_ready;                                                                      // rsp_xbar_mux_004:sink2_ready -> rsp_xbar_demux_016:src2_ready
	wire         rsp_xbar_demux_016_src3_endofpacket;                                                                // rsp_xbar_demux_016:src3_endofpacket -> rsp_xbar_mux_011:sink15_endofpacket
	wire         rsp_xbar_demux_016_src3_valid;                                                                      // rsp_xbar_demux_016:src3_valid -> rsp_xbar_mux_011:sink15_valid
	wire         rsp_xbar_demux_016_src3_startofpacket;                                                              // rsp_xbar_demux_016:src3_startofpacket -> rsp_xbar_mux_011:sink15_startofpacket
	wire  [94:0] rsp_xbar_demux_016_src3_data;                                                                       // rsp_xbar_demux_016:src3_data -> rsp_xbar_mux_011:sink15_data
	wire  [65:0] rsp_xbar_demux_016_src3_channel;                                                                    // rsp_xbar_demux_016:src3_channel -> rsp_xbar_mux_011:sink15_channel
	wire         rsp_xbar_demux_016_src3_ready;                                                                      // rsp_xbar_mux_011:sink15_ready -> rsp_xbar_demux_016:src3_ready
	wire         rsp_xbar_demux_017_src0_endofpacket;                                                                // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux:sink17_endofpacket
	wire         rsp_xbar_demux_017_src0_valid;                                                                      // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux:sink17_valid
	wire         rsp_xbar_demux_017_src0_startofpacket;                                                              // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux:sink17_startofpacket
	wire  [94:0] rsp_xbar_demux_017_src0_data;                                                                       // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux:sink17_data
	wire  [65:0] rsp_xbar_demux_017_src0_channel;                                                                    // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux:sink17_channel
	wire         rsp_xbar_demux_017_src0_ready;                                                                      // rsp_xbar_mux:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire         rsp_xbar_demux_017_src1_endofpacket;                                                                // rsp_xbar_demux_017:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_017_src1_valid;                                                                      // rsp_xbar_demux_017:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_017_src1_startofpacket;                                                              // rsp_xbar_demux_017:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_017_src1_data;                                                                       // rsp_xbar_demux_017:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [65:0] rsp_xbar_demux_017_src1_channel;                                                                    // rsp_xbar_demux_017:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_017_src1_ready;                                                                      // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux_017:src1_ready
	wire         rsp_xbar_demux_017_src2_endofpacket;                                                                // rsp_xbar_demux_017:src2_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire         rsp_xbar_demux_017_src2_valid;                                                                      // rsp_xbar_demux_017:src2_valid -> rsp_xbar_mux_002:sink0_valid
	wire         rsp_xbar_demux_017_src2_startofpacket;                                                              // rsp_xbar_demux_017:src2_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_017_src2_data;                                                                       // rsp_xbar_demux_017:src2_data -> rsp_xbar_mux_002:sink0_data
	wire  [65:0] rsp_xbar_demux_017_src2_channel;                                                                    // rsp_xbar_demux_017:src2_channel -> rsp_xbar_mux_002:sink0_channel
	wire         rsp_xbar_demux_017_src2_ready;                                                                      // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_017:src2_ready
	wire         rsp_xbar_demux_017_src3_endofpacket;                                                                // rsp_xbar_demux_017:src3_endofpacket -> rsp_xbar_mux_011:sink16_endofpacket
	wire         rsp_xbar_demux_017_src3_valid;                                                                      // rsp_xbar_demux_017:src3_valid -> rsp_xbar_mux_011:sink16_valid
	wire         rsp_xbar_demux_017_src3_startofpacket;                                                              // rsp_xbar_demux_017:src3_startofpacket -> rsp_xbar_mux_011:sink16_startofpacket
	wire  [94:0] rsp_xbar_demux_017_src3_data;                                                                       // rsp_xbar_demux_017:src3_data -> rsp_xbar_mux_011:sink16_data
	wire  [65:0] rsp_xbar_demux_017_src3_channel;                                                                    // rsp_xbar_demux_017:src3_channel -> rsp_xbar_mux_011:sink16_channel
	wire         rsp_xbar_demux_017_src3_ready;                                                                      // rsp_xbar_mux_011:sink16_ready -> rsp_xbar_demux_017:src3_ready
	wire         rsp_xbar_demux_018_src0_endofpacket;                                                                // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux:sink18_endofpacket
	wire         rsp_xbar_demux_018_src0_valid;                                                                      // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux:sink18_valid
	wire         rsp_xbar_demux_018_src0_startofpacket;                                                              // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux:sink18_startofpacket
	wire  [94:0] rsp_xbar_demux_018_src0_data;                                                                       // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux:sink18_data
	wire  [65:0] rsp_xbar_demux_018_src0_channel;                                                                    // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux:sink18_channel
	wire         rsp_xbar_demux_018_src0_ready;                                                                      // rsp_xbar_mux:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire         rsp_xbar_demux_018_src1_endofpacket;                                                                // rsp_xbar_demux_018:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_018_src1_valid;                                                                      // rsp_xbar_demux_018:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_018_src1_startofpacket;                                                              // rsp_xbar_demux_018:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_018_src1_data;                                                                       // rsp_xbar_demux_018:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [65:0] rsp_xbar_demux_018_src1_channel;                                                                    // rsp_xbar_demux_018:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_018_src1_ready;                                                                      // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_018:src1_ready
	wire         rsp_xbar_demux_018_src2_endofpacket;                                                                // rsp_xbar_demux_018:src2_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire         rsp_xbar_demux_018_src2_valid;                                                                      // rsp_xbar_demux_018:src2_valid -> rsp_xbar_mux_002:sink1_valid
	wire         rsp_xbar_demux_018_src2_startofpacket;                                                              // rsp_xbar_demux_018:src2_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_018_src2_data;                                                                       // rsp_xbar_demux_018:src2_data -> rsp_xbar_mux_002:sink1_data
	wire  [65:0] rsp_xbar_demux_018_src2_channel;                                                                    // rsp_xbar_demux_018:src2_channel -> rsp_xbar_mux_002:sink1_channel
	wire         rsp_xbar_demux_018_src2_ready;                                                                      // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_018:src2_ready
	wire         rsp_xbar_demux_018_src3_endofpacket;                                                                // rsp_xbar_demux_018:src3_endofpacket -> rsp_xbar_mux_011:sink17_endofpacket
	wire         rsp_xbar_demux_018_src3_valid;                                                                      // rsp_xbar_demux_018:src3_valid -> rsp_xbar_mux_011:sink17_valid
	wire         rsp_xbar_demux_018_src3_startofpacket;                                                              // rsp_xbar_demux_018:src3_startofpacket -> rsp_xbar_mux_011:sink17_startofpacket
	wire  [94:0] rsp_xbar_demux_018_src3_data;                                                                       // rsp_xbar_demux_018:src3_data -> rsp_xbar_mux_011:sink17_data
	wire  [65:0] rsp_xbar_demux_018_src3_channel;                                                                    // rsp_xbar_demux_018:src3_channel -> rsp_xbar_mux_011:sink17_channel
	wire         rsp_xbar_demux_018_src3_ready;                                                                      // rsp_xbar_mux_011:sink17_ready -> rsp_xbar_demux_018:src3_ready
	wire         rsp_xbar_demux_019_src0_endofpacket;                                                                // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux:sink19_endofpacket
	wire         rsp_xbar_demux_019_src0_valid;                                                                      // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux:sink19_valid
	wire         rsp_xbar_demux_019_src0_startofpacket;                                                              // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux:sink19_startofpacket
	wire  [94:0] rsp_xbar_demux_019_src0_data;                                                                       // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux:sink19_data
	wire  [65:0] rsp_xbar_demux_019_src0_channel;                                                                    // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux:sink19_channel
	wire         rsp_xbar_demux_019_src0_ready;                                                                      // rsp_xbar_mux:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire         rsp_xbar_demux_019_src1_endofpacket;                                                                // rsp_xbar_demux_019:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_019_src1_valid;                                                                      // rsp_xbar_demux_019:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_019_src1_startofpacket;                                                              // rsp_xbar_demux_019:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_019_src1_data;                                                                       // rsp_xbar_demux_019:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [65:0] rsp_xbar_demux_019_src1_channel;                                                                    // rsp_xbar_demux_019:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_019_src1_ready;                                                                      // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_019:src1_ready
	wire         rsp_xbar_demux_019_src2_endofpacket;                                                                // rsp_xbar_demux_019:src2_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire         rsp_xbar_demux_019_src2_valid;                                                                      // rsp_xbar_demux_019:src2_valid -> rsp_xbar_mux_002:sink2_valid
	wire         rsp_xbar_demux_019_src2_startofpacket;                                                              // rsp_xbar_demux_019:src2_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_019_src2_data;                                                                       // rsp_xbar_demux_019:src2_data -> rsp_xbar_mux_002:sink2_data
	wire  [65:0] rsp_xbar_demux_019_src2_channel;                                                                    // rsp_xbar_demux_019:src2_channel -> rsp_xbar_mux_002:sink2_channel
	wire         rsp_xbar_demux_019_src2_ready;                                                                      // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_019:src2_ready
	wire         rsp_xbar_demux_019_src3_endofpacket;                                                                // rsp_xbar_demux_019:src3_endofpacket -> rsp_xbar_mux_011:sink18_endofpacket
	wire         rsp_xbar_demux_019_src3_valid;                                                                      // rsp_xbar_demux_019:src3_valid -> rsp_xbar_mux_011:sink18_valid
	wire         rsp_xbar_demux_019_src3_startofpacket;                                                              // rsp_xbar_demux_019:src3_startofpacket -> rsp_xbar_mux_011:sink18_startofpacket
	wire  [94:0] rsp_xbar_demux_019_src3_data;                                                                       // rsp_xbar_demux_019:src3_data -> rsp_xbar_mux_011:sink18_data
	wire  [65:0] rsp_xbar_demux_019_src3_channel;                                                                    // rsp_xbar_demux_019:src3_channel -> rsp_xbar_mux_011:sink18_channel
	wire         rsp_xbar_demux_019_src3_ready;                                                                      // rsp_xbar_mux_011:sink18_ready -> rsp_xbar_demux_019:src3_ready
	wire         rsp_xbar_demux_020_src0_endofpacket;                                                                // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_020_src0_valid;                                                                      // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_020_src0_startofpacket;                                                              // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_020_src0_data;                                                                       // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink3_data
	wire  [65:0] rsp_xbar_demux_020_src0_channel;                                                                    // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_020_src0_ready;                                                                      // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_020:src0_ready
	wire         rsp_xbar_demux_021_src0_endofpacket;                                                                // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_021_src0_valid;                                                                      // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_021_src0_startofpacket;                                                              // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_021_src0_data;                                                                       // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink4_data
	wire  [65:0] rsp_xbar_demux_021_src0_channel;                                                                    // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_021_src0_ready;                                                                      // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_021:src0_ready
	wire         rsp_xbar_demux_021_src1_endofpacket;                                                                // rsp_xbar_demux_021:src1_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire         rsp_xbar_demux_021_src1_valid;                                                                      // rsp_xbar_demux_021:src1_valid -> rsp_xbar_mux_002:sink3_valid
	wire         rsp_xbar_demux_021_src1_startofpacket;                                                              // rsp_xbar_demux_021:src1_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_021_src1_data;                                                                       // rsp_xbar_demux_021:src1_data -> rsp_xbar_mux_002:sink3_data
	wire  [65:0] rsp_xbar_demux_021_src1_channel;                                                                    // rsp_xbar_demux_021:src1_channel -> rsp_xbar_mux_002:sink3_channel
	wire         rsp_xbar_demux_021_src1_ready;                                                                      // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_021:src1_ready
	wire         rsp_xbar_demux_022_src0_endofpacket;                                                                // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_022_src0_valid;                                                                      // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_022_src0_startofpacket;                                                              // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_022_src0_data;                                                                       // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [65:0] rsp_xbar_demux_022_src0_channel;                                                                    // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_022_src0_ready;                                                                      // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_022:src0_ready
	wire         rsp_xbar_demux_022_src1_endofpacket;                                                                // rsp_xbar_demux_022:src1_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	wire         rsp_xbar_demux_022_src1_valid;                                                                      // rsp_xbar_demux_022:src1_valid -> rsp_xbar_mux_002:sink4_valid
	wire         rsp_xbar_demux_022_src1_startofpacket;                                                              // rsp_xbar_demux_022:src1_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_022_src1_data;                                                                       // rsp_xbar_demux_022:src1_data -> rsp_xbar_mux_002:sink4_data
	wire  [65:0] rsp_xbar_demux_022_src1_channel;                                                                    // rsp_xbar_demux_022:src1_channel -> rsp_xbar_mux_002:sink4_channel
	wire         rsp_xbar_demux_022_src1_ready;                                                                      // rsp_xbar_mux_002:sink4_ready -> rsp_xbar_demux_022:src1_ready
	wire         rsp_xbar_demux_022_src2_endofpacket;                                                                // rsp_xbar_demux_022:src2_endofpacket -> rsp_xbar_mux_003:sink3_endofpacket
	wire         rsp_xbar_demux_022_src2_valid;                                                                      // rsp_xbar_demux_022:src2_valid -> rsp_xbar_mux_003:sink3_valid
	wire         rsp_xbar_demux_022_src2_startofpacket;                                                              // rsp_xbar_demux_022:src2_startofpacket -> rsp_xbar_mux_003:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_022_src2_data;                                                                       // rsp_xbar_demux_022:src2_data -> rsp_xbar_mux_003:sink3_data
	wire  [65:0] rsp_xbar_demux_022_src2_channel;                                                                    // rsp_xbar_demux_022:src2_channel -> rsp_xbar_mux_003:sink3_channel
	wire         rsp_xbar_demux_022_src2_ready;                                                                      // rsp_xbar_mux_003:sink3_ready -> rsp_xbar_demux_022:src2_ready
	wire         rsp_xbar_demux_022_src3_endofpacket;                                                                // rsp_xbar_demux_022:src3_endofpacket -> rsp_xbar_mux_004:sink3_endofpacket
	wire         rsp_xbar_demux_022_src3_valid;                                                                      // rsp_xbar_demux_022:src3_valid -> rsp_xbar_mux_004:sink3_valid
	wire         rsp_xbar_demux_022_src3_startofpacket;                                                              // rsp_xbar_demux_022:src3_startofpacket -> rsp_xbar_mux_004:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_022_src3_data;                                                                       // rsp_xbar_demux_022:src3_data -> rsp_xbar_mux_004:sink3_data
	wire  [65:0] rsp_xbar_demux_022_src3_channel;                                                                    // rsp_xbar_demux_022:src3_channel -> rsp_xbar_mux_004:sink3_channel
	wire         rsp_xbar_demux_022_src3_ready;                                                                      // rsp_xbar_mux_004:sink3_ready -> rsp_xbar_demux_022:src3_ready
	wire         rsp_xbar_demux_023_src0_endofpacket;                                                                // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_023_src0_valid;                                                                      // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_023_src0_startofpacket;                                                              // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_023_src0_data;                                                                       // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [65:0] rsp_xbar_demux_023_src0_channel;                                                                    // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_023_src0_ready;                                                                      // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_023:src0_ready
	wire         rsp_xbar_demux_023_src1_endofpacket;                                                                // rsp_xbar_demux_023:src1_endofpacket -> rsp_xbar_mux_002:sink5_endofpacket
	wire         rsp_xbar_demux_023_src1_valid;                                                                      // rsp_xbar_demux_023:src1_valid -> rsp_xbar_mux_002:sink5_valid
	wire         rsp_xbar_demux_023_src1_startofpacket;                                                              // rsp_xbar_demux_023:src1_startofpacket -> rsp_xbar_mux_002:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_023_src1_data;                                                                       // rsp_xbar_demux_023:src1_data -> rsp_xbar_mux_002:sink5_data
	wire  [65:0] rsp_xbar_demux_023_src1_channel;                                                                    // rsp_xbar_demux_023:src1_channel -> rsp_xbar_mux_002:sink5_channel
	wire         rsp_xbar_demux_023_src1_ready;                                                                      // rsp_xbar_mux_002:sink5_ready -> rsp_xbar_demux_023:src1_ready
	wire         rsp_xbar_demux_023_src2_endofpacket;                                                                // rsp_xbar_demux_023:src2_endofpacket -> rsp_xbar_mux_003:sink4_endofpacket
	wire         rsp_xbar_demux_023_src2_valid;                                                                      // rsp_xbar_demux_023:src2_valid -> rsp_xbar_mux_003:sink4_valid
	wire         rsp_xbar_demux_023_src2_startofpacket;                                                              // rsp_xbar_demux_023:src2_startofpacket -> rsp_xbar_mux_003:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_023_src2_data;                                                                       // rsp_xbar_demux_023:src2_data -> rsp_xbar_mux_003:sink4_data
	wire  [65:0] rsp_xbar_demux_023_src2_channel;                                                                    // rsp_xbar_demux_023:src2_channel -> rsp_xbar_mux_003:sink4_channel
	wire         rsp_xbar_demux_023_src2_ready;                                                                      // rsp_xbar_mux_003:sink4_ready -> rsp_xbar_demux_023:src2_ready
	wire         rsp_xbar_demux_023_src3_endofpacket;                                                                // rsp_xbar_demux_023:src3_endofpacket -> rsp_xbar_mux_004:sink4_endofpacket
	wire         rsp_xbar_demux_023_src3_valid;                                                                      // rsp_xbar_demux_023:src3_valid -> rsp_xbar_mux_004:sink4_valid
	wire         rsp_xbar_demux_023_src3_startofpacket;                                                              // rsp_xbar_demux_023:src3_startofpacket -> rsp_xbar_mux_004:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_023_src3_data;                                                                       // rsp_xbar_demux_023:src3_data -> rsp_xbar_mux_004:sink4_data
	wire  [65:0] rsp_xbar_demux_023_src3_channel;                                                                    // rsp_xbar_demux_023:src3_channel -> rsp_xbar_mux_004:sink4_channel
	wire         rsp_xbar_demux_023_src3_ready;                                                                      // rsp_xbar_mux_004:sink4_ready -> rsp_xbar_demux_023:src3_ready
	wire         rsp_xbar_demux_024_src0_endofpacket;                                                                // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_024_src0_valid;                                                                      // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_024_src0_startofpacket;                                                              // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_024_src0_data;                                                                       // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [65:0] rsp_xbar_demux_024_src0_channel;                                                                    // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_024_src0_ready;                                                                      // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_024:src0_ready
	wire         rsp_xbar_demux_024_src1_endofpacket;                                                                // rsp_xbar_demux_024:src1_endofpacket -> rsp_xbar_mux_002:sink6_endofpacket
	wire         rsp_xbar_demux_024_src1_valid;                                                                      // rsp_xbar_demux_024:src1_valid -> rsp_xbar_mux_002:sink6_valid
	wire         rsp_xbar_demux_024_src1_startofpacket;                                                              // rsp_xbar_demux_024:src1_startofpacket -> rsp_xbar_mux_002:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_024_src1_data;                                                                       // rsp_xbar_demux_024:src1_data -> rsp_xbar_mux_002:sink6_data
	wire  [65:0] rsp_xbar_demux_024_src1_channel;                                                                    // rsp_xbar_demux_024:src1_channel -> rsp_xbar_mux_002:sink6_channel
	wire         rsp_xbar_demux_024_src1_ready;                                                                      // rsp_xbar_mux_002:sink6_ready -> rsp_xbar_demux_024:src1_ready
	wire         rsp_xbar_demux_024_src2_endofpacket;                                                                // rsp_xbar_demux_024:src2_endofpacket -> rsp_xbar_mux_003:sink5_endofpacket
	wire         rsp_xbar_demux_024_src2_valid;                                                                      // rsp_xbar_demux_024:src2_valid -> rsp_xbar_mux_003:sink5_valid
	wire         rsp_xbar_demux_024_src2_startofpacket;                                                              // rsp_xbar_demux_024:src2_startofpacket -> rsp_xbar_mux_003:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_024_src2_data;                                                                       // rsp_xbar_demux_024:src2_data -> rsp_xbar_mux_003:sink5_data
	wire  [65:0] rsp_xbar_demux_024_src2_channel;                                                                    // rsp_xbar_demux_024:src2_channel -> rsp_xbar_mux_003:sink5_channel
	wire         rsp_xbar_demux_024_src2_ready;                                                                      // rsp_xbar_mux_003:sink5_ready -> rsp_xbar_demux_024:src2_ready
	wire         rsp_xbar_demux_024_src3_endofpacket;                                                                // rsp_xbar_demux_024:src3_endofpacket -> rsp_xbar_mux_004:sink5_endofpacket
	wire         rsp_xbar_demux_024_src3_valid;                                                                      // rsp_xbar_demux_024:src3_valid -> rsp_xbar_mux_004:sink5_valid
	wire         rsp_xbar_demux_024_src3_startofpacket;                                                              // rsp_xbar_demux_024:src3_startofpacket -> rsp_xbar_mux_004:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_024_src3_data;                                                                       // rsp_xbar_demux_024:src3_data -> rsp_xbar_mux_004:sink5_data
	wire  [65:0] rsp_xbar_demux_024_src3_channel;                                                                    // rsp_xbar_demux_024:src3_channel -> rsp_xbar_mux_004:sink5_channel
	wire         rsp_xbar_demux_024_src3_ready;                                                                      // rsp_xbar_mux_004:sink5_ready -> rsp_xbar_demux_024:src3_ready
	wire         rsp_xbar_demux_025_src0_endofpacket;                                                                // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_002:sink7_endofpacket
	wire         rsp_xbar_demux_025_src0_valid;                                                                      // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_002:sink7_valid
	wire         rsp_xbar_demux_025_src0_startofpacket;                                                              // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_002:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_025_src0_data;                                                                       // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_002:sink7_data
	wire  [65:0] rsp_xbar_demux_025_src0_channel;                                                                    // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_002:sink7_channel
	wire         rsp_xbar_demux_025_src0_ready;                                                                      // rsp_xbar_mux_002:sink7_ready -> rsp_xbar_demux_025:src0_ready
	wire         rsp_xbar_demux_026_src0_endofpacket;                                                                // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_002:sink8_endofpacket
	wire         rsp_xbar_demux_026_src0_valid;                                                                      // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_002:sink8_valid
	wire         rsp_xbar_demux_026_src0_startofpacket;                                                              // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_002:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_026_src0_data;                                                                       // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_002:sink8_data
	wire  [65:0] rsp_xbar_demux_026_src0_channel;                                                                    // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_002:sink8_channel
	wire         rsp_xbar_demux_026_src0_ready;                                                                      // rsp_xbar_mux_002:sink8_ready -> rsp_xbar_demux_026:src0_ready
	wire         rsp_xbar_demux_027_src0_endofpacket;                                                                // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_002:sink9_endofpacket
	wire         rsp_xbar_demux_027_src0_valid;                                                                      // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_002:sink9_valid
	wire         rsp_xbar_demux_027_src0_startofpacket;                                                              // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_002:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_027_src0_data;                                                                       // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_002:sink9_data
	wire  [65:0] rsp_xbar_demux_027_src0_channel;                                                                    // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_002:sink9_channel
	wire         rsp_xbar_demux_027_src0_ready;                                                                      // rsp_xbar_mux_002:sink9_ready -> rsp_xbar_demux_027:src0_ready
	wire         rsp_xbar_demux_028_src0_endofpacket;                                                                // rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux_002:sink10_endofpacket
	wire         rsp_xbar_demux_028_src0_valid;                                                                      // rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux_002:sink10_valid
	wire         rsp_xbar_demux_028_src0_startofpacket;                                                              // rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux_002:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_028_src0_data;                                                                       // rsp_xbar_demux_028:src0_data -> rsp_xbar_mux_002:sink10_data
	wire  [65:0] rsp_xbar_demux_028_src0_channel;                                                                    // rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux_002:sink10_channel
	wire         rsp_xbar_demux_028_src0_ready;                                                                      // rsp_xbar_mux_002:sink10_ready -> rsp_xbar_demux_028:src0_ready
	wire         rsp_xbar_demux_029_src0_endofpacket;                                                                // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_003:sink6_endofpacket
	wire         rsp_xbar_demux_029_src0_valid;                                                                      // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_003:sink6_valid
	wire         rsp_xbar_demux_029_src0_startofpacket;                                                              // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_003:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_029_src0_data;                                                                       // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_003:sink6_data
	wire  [65:0] rsp_xbar_demux_029_src0_channel;                                                                    // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_003:sink6_channel
	wire         rsp_xbar_demux_029_src0_ready;                                                                      // rsp_xbar_mux_003:sink6_ready -> rsp_xbar_demux_029:src0_ready
	wire         rsp_xbar_demux_030_src0_endofpacket;                                                                // rsp_xbar_demux_030:src0_endofpacket -> rsp_xbar_mux_003:sink7_endofpacket
	wire         rsp_xbar_demux_030_src0_valid;                                                                      // rsp_xbar_demux_030:src0_valid -> rsp_xbar_mux_003:sink7_valid
	wire         rsp_xbar_demux_030_src0_startofpacket;                                                              // rsp_xbar_demux_030:src0_startofpacket -> rsp_xbar_mux_003:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_030_src0_data;                                                                       // rsp_xbar_demux_030:src0_data -> rsp_xbar_mux_003:sink7_data
	wire  [65:0] rsp_xbar_demux_030_src0_channel;                                                                    // rsp_xbar_demux_030:src0_channel -> rsp_xbar_mux_003:sink7_channel
	wire         rsp_xbar_demux_030_src0_ready;                                                                      // rsp_xbar_mux_003:sink7_ready -> rsp_xbar_demux_030:src0_ready
	wire         rsp_xbar_demux_030_src1_endofpacket;                                                                // rsp_xbar_demux_030:src1_endofpacket -> rsp_xbar_mux_004:sink6_endofpacket
	wire         rsp_xbar_demux_030_src1_valid;                                                                      // rsp_xbar_demux_030:src1_valid -> rsp_xbar_mux_004:sink6_valid
	wire         rsp_xbar_demux_030_src1_startofpacket;                                                              // rsp_xbar_demux_030:src1_startofpacket -> rsp_xbar_mux_004:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_030_src1_data;                                                                       // rsp_xbar_demux_030:src1_data -> rsp_xbar_mux_004:sink6_data
	wire  [65:0] rsp_xbar_demux_030_src1_channel;                                                                    // rsp_xbar_demux_030:src1_channel -> rsp_xbar_mux_004:sink6_channel
	wire         rsp_xbar_demux_030_src1_ready;                                                                      // rsp_xbar_mux_004:sink6_ready -> rsp_xbar_demux_030:src1_ready
	wire         rsp_xbar_demux_031_src0_endofpacket;                                                                // rsp_xbar_demux_031:src0_endofpacket -> rsp_xbar_mux_003:sink8_endofpacket
	wire         rsp_xbar_demux_031_src0_valid;                                                                      // rsp_xbar_demux_031:src0_valid -> rsp_xbar_mux_003:sink8_valid
	wire         rsp_xbar_demux_031_src0_startofpacket;                                                              // rsp_xbar_demux_031:src0_startofpacket -> rsp_xbar_mux_003:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_031_src0_data;                                                                       // rsp_xbar_demux_031:src0_data -> rsp_xbar_mux_003:sink8_data
	wire  [65:0] rsp_xbar_demux_031_src0_channel;                                                                    // rsp_xbar_demux_031:src0_channel -> rsp_xbar_mux_003:sink8_channel
	wire         rsp_xbar_demux_031_src0_ready;                                                                      // rsp_xbar_mux_003:sink8_ready -> rsp_xbar_demux_031:src0_ready
	wire         rsp_xbar_demux_031_src1_endofpacket;                                                                // rsp_xbar_demux_031:src1_endofpacket -> rsp_xbar_mux_004:sink7_endofpacket
	wire         rsp_xbar_demux_031_src1_valid;                                                                      // rsp_xbar_demux_031:src1_valid -> rsp_xbar_mux_004:sink7_valid
	wire         rsp_xbar_demux_031_src1_startofpacket;                                                              // rsp_xbar_demux_031:src1_startofpacket -> rsp_xbar_mux_004:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_031_src1_data;                                                                       // rsp_xbar_demux_031:src1_data -> rsp_xbar_mux_004:sink7_data
	wire  [65:0] rsp_xbar_demux_031_src1_channel;                                                                    // rsp_xbar_demux_031:src1_channel -> rsp_xbar_mux_004:sink7_channel
	wire         rsp_xbar_demux_031_src1_ready;                                                                      // rsp_xbar_mux_004:sink7_ready -> rsp_xbar_demux_031:src1_ready
	wire         rsp_xbar_demux_031_src2_endofpacket;                                                                // rsp_xbar_demux_031:src2_endofpacket -> rsp_xbar_mux_005:sink3_endofpacket
	wire         rsp_xbar_demux_031_src2_valid;                                                                      // rsp_xbar_demux_031:src2_valid -> rsp_xbar_mux_005:sink3_valid
	wire         rsp_xbar_demux_031_src2_startofpacket;                                                              // rsp_xbar_demux_031:src2_startofpacket -> rsp_xbar_mux_005:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_031_src2_data;                                                                       // rsp_xbar_demux_031:src2_data -> rsp_xbar_mux_005:sink3_data
	wire  [65:0] rsp_xbar_demux_031_src2_channel;                                                                    // rsp_xbar_demux_031:src2_channel -> rsp_xbar_mux_005:sink3_channel
	wire         rsp_xbar_demux_031_src2_ready;                                                                      // rsp_xbar_mux_005:sink3_ready -> rsp_xbar_demux_031:src2_ready
	wire         rsp_xbar_demux_031_src3_endofpacket;                                                                // rsp_xbar_demux_031:src3_endofpacket -> rsp_xbar_mux_006:sink3_endofpacket
	wire         rsp_xbar_demux_031_src3_valid;                                                                      // rsp_xbar_demux_031:src3_valid -> rsp_xbar_mux_006:sink3_valid
	wire         rsp_xbar_demux_031_src3_startofpacket;                                                              // rsp_xbar_demux_031:src3_startofpacket -> rsp_xbar_mux_006:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_031_src3_data;                                                                       // rsp_xbar_demux_031:src3_data -> rsp_xbar_mux_006:sink3_data
	wire  [65:0] rsp_xbar_demux_031_src3_channel;                                                                    // rsp_xbar_demux_031:src3_channel -> rsp_xbar_mux_006:sink3_channel
	wire         rsp_xbar_demux_031_src3_ready;                                                                      // rsp_xbar_mux_006:sink3_ready -> rsp_xbar_demux_031:src3_ready
	wire         rsp_xbar_demux_032_src0_endofpacket;                                                                // rsp_xbar_demux_032:src0_endofpacket -> rsp_xbar_mux_003:sink9_endofpacket
	wire         rsp_xbar_demux_032_src0_valid;                                                                      // rsp_xbar_demux_032:src0_valid -> rsp_xbar_mux_003:sink9_valid
	wire         rsp_xbar_demux_032_src0_startofpacket;                                                              // rsp_xbar_demux_032:src0_startofpacket -> rsp_xbar_mux_003:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_032_src0_data;                                                                       // rsp_xbar_demux_032:src0_data -> rsp_xbar_mux_003:sink9_data
	wire  [65:0] rsp_xbar_demux_032_src0_channel;                                                                    // rsp_xbar_demux_032:src0_channel -> rsp_xbar_mux_003:sink9_channel
	wire         rsp_xbar_demux_032_src0_ready;                                                                      // rsp_xbar_mux_003:sink9_ready -> rsp_xbar_demux_032:src0_ready
	wire         rsp_xbar_demux_032_src1_endofpacket;                                                                // rsp_xbar_demux_032:src1_endofpacket -> rsp_xbar_mux_004:sink8_endofpacket
	wire         rsp_xbar_demux_032_src1_valid;                                                                      // rsp_xbar_demux_032:src1_valid -> rsp_xbar_mux_004:sink8_valid
	wire         rsp_xbar_demux_032_src1_startofpacket;                                                              // rsp_xbar_demux_032:src1_startofpacket -> rsp_xbar_mux_004:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_032_src1_data;                                                                       // rsp_xbar_demux_032:src1_data -> rsp_xbar_mux_004:sink8_data
	wire  [65:0] rsp_xbar_demux_032_src1_channel;                                                                    // rsp_xbar_demux_032:src1_channel -> rsp_xbar_mux_004:sink8_channel
	wire         rsp_xbar_demux_032_src1_ready;                                                                      // rsp_xbar_mux_004:sink8_ready -> rsp_xbar_demux_032:src1_ready
	wire         rsp_xbar_demux_032_src2_endofpacket;                                                                // rsp_xbar_demux_032:src2_endofpacket -> rsp_xbar_mux_005:sink4_endofpacket
	wire         rsp_xbar_demux_032_src2_valid;                                                                      // rsp_xbar_demux_032:src2_valid -> rsp_xbar_mux_005:sink4_valid
	wire         rsp_xbar_demux_032_src2_startofpacket;                                                              // rsp_xbar_demux_032:src2_startofpacket -> rsp_xbar_mux_005:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_032_src2_data;                                                                       // rsp_xbar_demux_032:src2_data -> rsp_xbar_mux_005:sink4_data
	wire  [65:0] rsp_xbar_demux_032_src2_channel;                                                                    // rsp_xbar_demux_032:src2_channel -> rsp_xbar_mux_005:sink4_channel
	wire         rsp_xbar_demux_032_src2_ready;                                                                      // rsp_xbar_mux_005:sink4_ready -> rsp_xbar_demux_032:src2_ready
	wire         rsp_xbar_demux_032_src3_endofpacket;                                                                // rsp_xbar_demux_032:src3_endofpacket -> rsp_xbar_mux_006:sink4_endofpacket
	wire         rsp_xbar_demux_032_src3_valid;                                                                      // rsp_xbar_demux_032:src3_valid -> rsp_xbar_mux_006:sink4_valid
	wire         rsp_xbar_demux_032_src3_startofpacket;                                                              // rsp_xbar_demux_032:src3_startofpacket -> rsp_xbar_mux_006:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_032_src3_data;                                                                       // rsp_xbar_demux_032:src3_data -> rsp_xbar_mux_006:sink4_data
	wire  [65:0] rsp_xbar_demux_032_src3_channel;                                                                    // rsp_xbar_demux_032:src3_channel -> rsp_xbar_mux_006:sink4_channel
	wire         rsp_xbar_demux_032_src3_ready;                                                                      // rsp_xbar_mux_006:sink4_ready -> rsp_xbar_demux_032:src3_ready
	wire         rsp_xbar_demux_033_src0_endofpacket;                                                                // rsp_xbar_demux_033:src0_endofpacket -> rsp_xbar_mux_003:sink10_endofpacket
	wire         rsp_xbar_demux_033_src0_valid;                                                                      // rsp_xbar_demux_033:src0_valid -> rsp_xbar_mux_003:sink10_valid
	wire         rsp_xbar_demux_033_src0_startofpacket;                                                              // rsp_xbar_demux_033:src0_startofpacket -> rsp_xbar_mux_003:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_033_src0_data;                                                                       // rsp_xbar_demux_033:src0_data -> rsp_xbar_mux_003:sink10_data
	wire  [65:0] rsp_xbar_demux_033_src0_channel;                                                                    // rsp_xbar_demux_033:src0_channel -> rsp_xbar_mux_003:sink10_channel
	wire         rsp_xbar_demux_033_src0_ready;                                                                      // rsp_xbar_mux_003:sink10_ready -> rsp_xbar_demux_033:src0_ready
	wire         rsp_xbar_demux_033_src1_endofpacket;                                                                // rsp_xbar_demux_033:src1_endofpacket -> rsp_xbar_mux_004:sink9_endofpacket
	wire         rsp_xbar_demux_033_src1_valid;                                                                      // rsp_xbar_demux_033:src1_valid -> rsp_xbar_mux_004:sink9_valid
	wire         rsp_xbar_demux_033_src1_startofpacket;                                                              // rsp_xbar_demux_033:src1_startofpacket -> rsp_xbar_mux_004:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_033_src1_data;                                                                       // rsp_xbar_demux_033:src1_data -> rsp_xbar_mux_004:sink9_data
	wire  [65:0] rsp_xbar_demux_033_src1_channel;                                                                    // rsp_xbar_demux_033:src1_channel -> rsp_xbar_mux_004:sink9_channel
	wire         rsp_xbar_demux_033_src1_ready;                                                                      // rsp_xbar_mux_004:sink9_ready -> rsp_xbar_demux_033:src1_ready
	wire         rsp_xbar_demux_033_src2_endofpacket;                                                                // rsp_xbar_demux_033:src2_endofpacket -> rsp_xbar_mux_005:sink5_endofpacket
	wire         rsp_xbar_demux_033_src2_valid;                                                                      // rsp_xbar_demux_033:src2_valid -> rsp_xbar_mux_005:sink5_valid
	wire         rsp_xbar_demux_033_src2_startofpacket;                                                              // rsp_xbar_demux_033:src2_startofpacket -> rsp_xbar_mux_005:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_033_src2_data;                                                                       // rsp_xbar_demux_033:src2_data -> rsp_xbar_mux_005:sink5_data
	wire  [65:0] rsp_xbar_demux_033_src2_channel;                                                                    // rsp_xbar_demux_033:src2_channel -> rsp_xbar_mux_005:sink5_channel
	wire         rsp_xbar_demux_033_src2_ready;                                                                      // rsp_xbar_mux_005:sink5_ready -> rsp_xbar_demux_033:src2_ready
	wire         rsp_xbar_demux_033_src3_endofpacket;                                                                // rsp_xbar_demux_033:src3_endofpacket -> rsp_xbar_mux_006:sink5_endofpacket
	wire         rsp_xbar_demux_033_src3_valid;                                                                      // rsp_xbar_demux_033:src3_valid -> rsp_xbar_mux_006:sink5_valid
	wire         rsp_xbar_demux_033_src3_startofpacket;                                                              // rsp_xbar_demux_033:src3_startofpacket -> rsp_xbar_mux_006:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_033_src3_data;                                                                       // rsp_xbar_demux_033:src3_data -> rsp_xbar_mux_006:sink5_data
	wire  [65:0] rsp_xbar_demux_033_src3_channel;                                                                    // rsp_xbar_demux_033:src3_channel -> rsp_xbar_mux_006:sink5_channel
	wire         rsp_xbar_demux_033_src3_ready;                                                                      // rsp_xbar_mux_006:sink5_ready -> rsp_xbar_demux_033:src3_ready
	wire         rsp_xbar_demux_034_src0_endofpacket;                                                                // rsp_xbar_demux_034:src0_endofpacket -> rsp_xbar_mux_004:sink10_endofpacket
	wire         rsp_xbar_demux_034_src0_valid;                                                                      // rsp_xbar_demux_034:src0_valid -> rsp_xbar_mux_004:sink10_valid
	wire         rsp_xbar_demux_034_src0_startofpacket;                                                              // rsp_xbar_demux_034:src0_startofpacket -> rsp_xbar_mux_004:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_034_src0_data;                                                                       // rsp_xbar_demux_034:src0_data -> rsp_xbar_mux_004:sink10_data
	wire  [65:0] rsp_xbar_demux_034_src0_channel;                                                                    // rsp_xbar_demux_034:src0_channel -> rsp_xbar_mux_004:sink10_channel
	wire         rsp_xbar_demux_034_src0_ready;                                                                      // rsp_xbar_mux_004:sink10_ready -> rsp_xbar_demux_034:src0_ready
	wire         rsp_xbar_demux_035_src0_endofpacket;                                                                // rsp_xbar_demux_035:src0_endofpacket -> rsp_xbar_mux_004:sink11_endofpacket
	wire         rsp_xbar_demux_035_src0_valid;                                                                      // rsp_xbar_demux_035:src0_valid -> rsp_xbar_mux_004:sink11_valid
	wire         rsp_xbar_demux_035_src0_startofpacket;                                                              // rsp_xbar_demux_035:src0_startofpacket -> rsp_xbar_mux_004:sink11_startofpacket
	wire  [94:0] rsp_xbar_demux_035_src0_data;                                                                       // rsp_xbar_demux_035:src0_data -> rsp_xbar_mux_004:sink11_data
	wire  [65:0] rsp_xbar_demux_035_src0_channel;                                                                    // rsp_xbar_demux_035:src0_channel -> rsp_xbar_mux_004:sink11_channel
	wire         rsp_xbar_demux_035_src0_ready;                                                                      // rsp_xbar_mux_004:sink11_ready -> rsp_xbar_demux_035:src0_ready
	wire         rsp_xbar_demux_036_src0_endofpacket;                                                                // rsp_xbar_demux_036:src0_endofpacket -> rsp_xbar_mux_004:sink12_endofpacket
	wire         rsp_xbar_demux_036_src0_valid;                                                                      // rsp_xbar_demux_036:src0_valid -> rsp_xbar_mux_004:sink12_valid
	wire         rsp_xbar_demux_036_src0_startofpacket;                                                              // rsp_xbar_demux_036:src0_startofpacket -> rsp_xbar_mux_004:sink12_startofpacket
	wire  [94:0] rsp_xbar_demux_036_src0_data;                                                                       // rsp_xbar_demux_036:src0_data -> rsp_xbar_mux_004:sink12_data
	wire  [65:0] rsp_xbar_demux_036_src0_channel;                                                                    // rsp_xbar_demux_036:src0_channel -> rsp_xbar_mux_004:sink12_channel
	wire         rsp_xbar_demux_036_src0_ready;                                                                      // rsp_xbar_mux_004:sink12_ready -> rsp_xbar_demux_036:src0_ready
	wire         rsp_xbar_demux_037_src0_endofpacket;                                                                // rsp_xbar_demux_037:src0_endofpacket -> rsp_xbar_mux_004:sink13_endofpacket
	wire         rsp_xbar_demux_037_src0_valid;                                                                      // rsp_xbar_demux_037:src0_valid -> rsp_xbar_mux_004:sink13_valid
	wire         rsp_xbar_demux_037_src0_startofpacket;                                                              // rsp_xbar_demux_037:src0_startofpacket -> rsp_xbar_mux_004:sink13_startofpacket
	wire  [94:0] rsp_xbar_demux_037_src0_data;                                                                       // rsp_xbar_demux_037:src0_data -> rsp_xbar_mux_004:sink13_data
	wire  [65:0] rsp_xbar_demux_037_src0_channel;                                                                    // rsp_xbar_demux_037:src0_channel -> rsp_xbar_mux_004:sink13_channel
	wire         rsp_xbar_demux_037_src0_ready;                                                                      // rsp_xbar_mux_004:sink13_ready -> rsp_xbar_demux_037:src0_ready
	wire         rsp_xbar_demux_038_src0_endofpacket;                                                                // rsp_xbar_demux_038:src0_endofpacket -> rsp_xbar_mux_005:sink6_endofpacket
	wire         rsp_xbar_demux_038_src0_valid;                                                                      // rsp_xbar_demux_038:src0_valid -> rsp_xbar_mux_005:sink6_valid
	wire         rsp_xbar_demux_038_src0_startofpacket;                                                              // rsp_xbar_demux_038:src0_startofpacket -> rsp_xbar_mux_005:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_038_src0_data;                                                                       // rsp_xbar_demux_038:src0_data -> rsp_xbar_mux_005:sink6_data
	wire  [65:0] rsp_xbar_demux_038_src0_channel;                                                                    // rsp_xbar_demux_038:src0_channel -> rsp_xbar_mux_005:sink6_channel
	wire         rsp_xbar_demux_038_src0_ready;                                                                      // rsp_xbar_mux_005:sink6_ready -> rsp_xbar_demux_038:src0_ready
	wire         rsp_xbar_demux_039_src0_endofpacket;                                                                // rsp_xbar_demux_039:src0_endofpacket -> rsp_xbar_mux_005:sink7_endofpacket
	wire         rsp_xbar_demux_039_src0_valid;                                                                      // rsp_xbar_demux_039:src0_valid -> rsp_xbar_mux_005:sink7_valid
	wire         rsp_xbar_demux_039_src0_startofpacket;                                                              // rsp_xbar_demux_039:src0_startofpacket -> rsp_xbar_mux_005:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_039_src0_data;                                                                       // rsp_xbar_demux_039:src0_data -> rsp_xbar_mux_005:sink7_data
	wire  [65:0] rsp_xbar_demux_039_src0_channel;                                                                    // rsp_xbar_demux_039:src0_channel -> rsp_xbar_mux_005:sink7_channel
	wire         rsp_xbar_demux_039_src0_ready;                                                                      // rsp_xbar_mux_005:sink7_ready -> rsp_xbar_demux_039:src0_ready
	wire         rsp_xbar_demux_039_src1_endofpacket;                                                                // rsp_xbar_demux_039:src1_endofpacket -> rsp_xbar_mux_006:sink6_endofpacket
	wire         rsp_xbar_demux_039_src1_valid;                                                                      // rsp_xbar_demux_039:src1_valid -> rsp_xbar_mux_006:sink6_valid
	wire         rsp_xbar_demux_039_src1_startofpacket;                                                              // rsp_xbar_demux_039:src1_startofpacket -> rsp_xbar_mux_006:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_039_src1_data;                                                                       // rsp_xbar_demux_039:src1_data -> rsp_xbar_mux_006:sink6_data
	wire  [65:0] rsp_xbar_demux_039_src1_channel;                                                                    // rsp_xbar_demux_039:src1_channel -> rsp_xbar_mux_006:sink6_channel
	wire         rsp_xbar_demux_039_src1_ready;                                                                      // rsp_xbar_mux_006:sink6_ready -> rsp_xbar_demux_039:src1_ready
	wire         rsp_xbar_demux_040_src0_endofpacket;                                                                // rsp_xbar_demux_040:src0_endofpacket -> rsp_xbar_mux_005:sink8_endofpacket
	wire         rsp_xbar_demux_040_src0_valid;                                                                      // rsp_xbar_demux_040:src0_valid -> rsp_xbar_mux_005:sink8_valid
	wire         rsp_xbar_demux_040_src0_startofpacket;                                                              // rsp_xbar_demux_040:src0_startofpacket -> rsp_xbar_mux_005:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_040_src0_data;                                                                       // rsp_xbar_demux_040:src0_data -> rsp_xbar_mux_005:sink8_data
	wire  [65:0] rsp_xbar_demux_040_src0_channel;                                                                    // rsp_xbar_demux_040:src0_channel -> rsp_xbar_mux_005:sink8_channel
	wire         rsp_xbar_demux_040_src0_ready;                                                                      // rsp_xbar_mux_005:sink8_ready -> rsp_xbar_demux_040:src0_ready
	wire         rsp_xbar_demux_040_src1_endofpacket;                                                                // rsp_xbar_demux_040:src1_endofpacket -> rsp_xbar_mux_006:sink7_endofpacket
	wire         rsp_xbar_demux_040_src1_valid;                                                                      // rsp_xbar_demux_040:src1_valid -> rsp_xbar_mux_006:sink7_valid
	wire         rsp_xbar_demux_040_src1_startofpacket;                                                              // rsp_xbar_demux_040:src1_startofpacket -> rsp_xbar_mux_006:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_040_src1_data;                                                                       // rsp_xbar_demux_040:src1_data -> rsp_xbar_mux_006:sink7_data
	wire  [65:0] rsp_xbar_demux_040_src1_channel;                                                                    // rsp_xbar_demux_040:src1_channel -> rsp_xbar_mux_006:sink7_channel
	wire         rsp_xbar_demux_040_src1_ready;                                                                      // rsp_xbar_mux_006:sink7_ready -> rsp_xbar_demux_040:src1_ready
	wire         rsp_xbar_demux_040_src2_endofpacket;                                                                // rsp_xbar_demux_040:src2_endofpacket -> rsp_xbar_mux_007:sink0_endofpacket
	wire         rsp_xbar_demux_040_src2_valid;                                                                      // rsp_xbar_demux_040:src2_valid -> rsp_xbar_mux_007:sink0_valid
	wire         rsp_xbar_demux_040_src2_startofpacket;                                                              // rsp_xbar_demux_040:src2_startofpacket -> rsp_xbar_mux_007:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_040_src2_data;                                                                       // rsp_xbar_demux_040:src2_data -> rsp_xbar_mux_007:sink0_data
	wire  [65:0] rsp_xbar_demux_040_src2_channel;                                                                    // rsp_xbar_demux_040:src2_channel -> rsp_xbar_mux_007:sink0_channel
	wire         rsp_xbar_demux_040_src2_ready;                                                                      // rsp_xbar_mux_007:sink0_ready -> rsp_xbar_demux_040:src2_ready
	wire         rsp_xbar_demux_040_src3_endofpacket;                                                                // rsp_xbar_demux_040:src3_endofpacket -> rsp_xbar_mux_008:sink0_endofpacket
	wire         rsp_xbar_demux_040_src3_valid;                                                                      // rsp_xbar_demux_040:src3_valid -> rsp_xbar_mux_008:sink0_valid
	wire         rsp_xbar_demux_040_src3_startofpacket;                                                              // rsp_xbar_demux_040:src3_startofpacket -> rsp_xbar_mux_008:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_040_src3_data;                                                                       // rsp_xbar_demux_040:src3_data -> rsp_xbar_mux_008:sink0_data
	wire  [65:0] rsp_xbar_demux_040_src3_channel;                                                                    // rsp_xbar_demux_040:src3_channel -> rsp_xbar_mux_008:sink0_channel
	wire         rsp_xbar_demux_040_src3_ready;                                                                      // rsp_xbar_mux_008:sink0_ready -> rsp_xbar_demux_040:src3_ready
	wire         rsp_xbar_demux_041_src0_endofpacket;                                                                // rsp_xbar_demux_041:src0_endofpacket -> rsp_xbar_mux_005:sink9_endofpacket
	wire         rsp_xbar_demux_041_src0_valid;                                                                      // rsp_xbar_demux_041:src0_valid -> rsp_xbar_mux_005:sink9_valid
	wire         rsp_xbar_demux_041_src0_startofpacket;                                                              // rsp_xbar_demux_041:src0_startofpacket -> rsp_xbar_mux_005:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_041_src0_data;                                                                       // rsp_xbar_demux_041:src0_data -> rsp_xbar_mux_005:sink9_data
	wire  [65:0] rsp_xbar_demux_041_src0_channel;                                                                    // rsp_xbar_demux_041:src0_channel -> rsp_xbar_mux_005:sink9_channel
	wire         rsp_xbar_demux_041_src0_ready;                                                                      // rsp_xbar_mux_005:sink9_ready -> rsp_xbar_demux_041:src0_ready
	wire         rsp_xbar_demux_041_src1_endofpacket;                                                                // rsp_xbar_demux_041:src1_endofpacket -> rsp_xbar_mux_006:sink8_endofpacket
	wire         rsp_xbar_demux_041_src1_valid;                                                                      // rsp_xbar_demux_041:src1_valid -> rsp_xbar_mux_006:sink8_valid
	wire         rsp_xbar_demux_041_src1_startofpacket;                                                              // rsp_xbar_demux_041:src1_startofpacket -> rsp_xbar_mux_006:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_041_src1_data;                                                                       // rsp_xbar_demux_041:src1_data -> rsp_xbar_mux_006:sink8_data
	wire  [65:0] rsp_xbar_demux_041_src1_channel;                                                                    // rsp_xbar_demux_041:src1_channel -> rsp_xbar_mux_006:sink8_channel
	wire         rsp_xbar_demux_041_src1_ready;                                                                      // rsp_xbar_mux_006:sink8_ready -> rsp_xbar_demux_041:src1_ready
	wire         rsp_xbar_demux_041_src2_endofpacket;                                                                // rsp_xbar_demux_041:src2_endofpacket -> rsp_xbar_mux_007:sink1_endofpacket
	wire         rsp_xbar_demux_041_src2_valid;                                                                      // rsp_xbar_demux_041:src2_valid -> rsp_xbar_mux_007:sink1_valid
	wire         rsp_xbar_demux_041_src2_startofpacket;                                                              // rsp_xbar_demux_041:src2_startofpacket -> rsp_xbar_mux_007:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_041_src2_data;                                                                       // rsp_xbar_demux_041:src2_data -> rsp_xbar_mux_007:sink1_data
	wire  [65:0] rsp_xbar_demux_041_src2_channel;                                                                    // rsp_xbar_demux_041:src2_channel -> rsp_xbar_mux_007:sink1_channel
	wire         rsp_xbar_demux_041_src2_ready;                                                                      // rsp_xbar_mux_007:sink1_ready -> rsp_xbar_demux_041:src2_ready
	wire         rsp_xbar_demux_041_src3_endofpacket;                                                                // rsp_xbar_demux_041:src3_endofpacket -> rsp_xbar_mux_008:sink1_endofpacket
	wire         rsp_xbar_demux_041_src3_valid;                                                                      // rsp_xbar_demux_041:src3_valid -> rsp_xbar_mux_008:sink1_valid
	wire         rsp_xbar_demux_041_src3_startofpacket;                                                              // rsp_xbar_demux_041:src3_startofpacket -> rsp_xbar_mux_008:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_041_src3_data;                                                                       // rsp_xbar_demux_041:src3_data -> rsp_xbar_mux_008:sink1_data
	wire  [65:0] rsp_xbar_demux_041_src3_channel;                                                                    // rsp_xbar_demux_041:src3_channel -> rsp_xbar_mux_008:sink1_channel
	wire         rsp_xbar_demux_041_src3_ready;                                                                      // rsp_xbar_mux_008:sink1_ready -> rsp_xbar_demux_041:src3_ready
	wire         rsp_xbar_demux_042_src0_endofpacket;                                                                // rsp_xbar_demux_042:src0_endofpacket -> rsp_xbar_mux_005:sink10_endofpacket
	wire         rsp_xbar_demux_042_src0_valid;                                                                      // rsp_xbar_demux_042:src0_valid -> rsp_xbar_mux_005:sink10_valid
	wire         rsp_xbar_demux_042_src0_startofpacket;                                                              // rsp_xbar_demux_042:src0_startofpacket -> rsp_xbar_mux_005:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_042_src0_data;                                                                       // rsp_xbar_demux_042:src0_data -> rsp_xbar_mux_005:sink10_data
	wire  [65:0] rsp_xbar_demux_042_src0_channel;                                                                    // rsp_xbar_demux_042:src0_channel -> rsp_xbar_mux_005:sink10_channel
	wire         rsp_xbar_demux_042_src0_ready;                                                                      // rsp_xbar_mux_005:sink10_ready -> rsp_xbar_demux_042:src0_ready
	wire         rsp_xbar_demux_042_src1_endofpacket;                                                                // rsp_xbar_demux_042:src1_endofpacket -> rsp_xbar_mux_006:sink9_endofpacket
	wire         rsp_xbar_demux_042_src1_valid;                                                                      // rsp_xbar_demux_042:src1_valid -> rsp_xbar_mux_006:sink9_valid
	wire         rsp_xbar_demux_042_src1_startofpacket;                                                              // rsp_xbar_demux_042:src1_startofpacket -> rsp_xbar_mux_006:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_042_src1_data;                                                                       // rsp_xbar_demux_042:src1_data -> rsp_xbar_mux_006:sink9_data
	wire  [65:0] rsp_xbar_demux_042_src1_channel;                                                                    // rsp_xbar_demux_042:src1_channel -> rsp_xbar_mux_006:sink9_channel
	wire         rsp_xbar_demux_042_src1_ready;                                                                      // rsp_xbar_mux_006:sink9_ready -> rsp_xbar_demux_042:src1_ready
	wire         rsp_xbar_demux_042_src2_endofpacket;                                                                // rsp_xbar_demux_042:src2_endofpacket -> rsp_xbar_mux_007:sink2_endofpacket
	wire         rsp_xbar_demux_042_src2_valid;                                                                      // rsp_xbar_demux_042:src2_valid -> rsp_xbar_mux_007:sink2_valid
	wire         rsp_xbar_demux_042_src2_startofpacket;                                                              // rsp_xbar_demux_042:src2_startofpacket -> rsp_xbar_mux_007:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_042_src2_data;                                                                       // rsp_xbar_demux_042:src2_data -> rsp_xbar_mux_007:sink2_data
	wire  [65:0] rsp_xbar_demux_042_src2_channel;                                                                    // rsp_xbar_demux_042:src2_channel -> rsp_xbar_mux_007:sink2_channel
	wire         rsp_xbar_demux_042_src2_ready;                                                                      // rsp_xbar_mux_007:sink2_ready -> rsp_xbar_demux_042:src2_ready
	wire         rsp_xbar_demux_042_src3_endofpacket;                                                                // rsp_xbar_demux_042:src3_endofpacket -> rsp_xbar_mux_008:sink2_endofpacket
	wire         rsp_xbar_demux_042_src3_valid;                                                                      // rsp_xbar_demux_042:src3_valid -> rsp_xbar_mux_008:sink2_valid
	wire         rsp_xbar_demux_042_src3_startofpacket;                                                              // rsp_xbar_demux_042:src3_startofpacket -> rsp_xbar_mux_008:sink2_startofpacket
	wire  [94:0] rsp_xbar_demux_042_src3_data;                                                                       // rsp_xbar_demux_042:src3_data -> rsp_xbar_mux_008:sink2_data
	wire  [65:0] rsp_xbar_demux_042_src3_channel;                                                                    // rsp_xbar_demux_042:src3_channel -> rsp_xbar_mux_008:sink2_channel
	wire         rsp_xbar_demux_042_src3_ready;                                                                      // rsp_xbar_mux_008:sink2_ready -> rsp_xbar_demux_042:src3_ready
	wire         rsp_xbar_demux_043_src0_endofpacket;                                                                // rsp_xbar_demux_043:src0_endofpacket -> rsp_xbar_mux_006:sink10_endofpacket
	wire         rsp_xbar_demux_043_src0_valid;                                                                      // rsp_xbar_demux_043:src0_valid -> rsp_xbar_mux_006:sink10_valid
	wire         rsp_xbar_demux_043_src0_startofpacket;                                                              // rsp_xbar_demux_043:src0_startofpacket -> rsp_xbar_mux_006:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_043_src0_data;                                                                       // rsp_xbar_demux_043:src0_data -> rsp_xbar_mux_006:sink10_data
	wire  [65:0] rsp_xbar_demux_043_src0_channel;                                                                    // rsp_xbar_demux_043:src0_channel -> rsp_xbar_mux_006:sink10_channel
	wire         rsp_xbar_demux_043_src0_ready;                                                                      // rsp_xbar_mux_006:sink10_ready -> rsp_xbar_demux_043:src0_ready
	wire         rsp_xbar_demux_044_src0_endofpacket;                                                                // rsp_xbar_demux_044:src0_endofpacket -> rsp_xbar_mux_006:sink11_endofpacket
	wire         rsp_xbar_demux_044_src0_valid;                                                                      // rsp_xbar_demux_044:src0_valid -> rsp_xbar_mux_006:sink11_valid
	wire         rsp_xbar_demux_044_src0_startofpacket;                                                              // rsp_xbar_demux_044:src0_startofpacket -> rsp_xbar_mux_006:sink11_startofpacket
	wire  [94:0] rsp_xbar_demux_044_src0_data;                                                                       // rsp_xbar_demux_044:src0_data -> rsp_xbar_mux_006:sink11_data
	wire  [65:0] rsp_xbar_demux_044_src0_channel;                                                                    // rsp_xbar_demux_044:src0_channel -> rsp_xbar_mux_006:sink11_channel
	wire         rsp_xbar_demux_044_src0_ready;                                                                      // rsp_xbar_mux_006:sink11_ready -> rsp_xbar_demux_044:src0_ready
	wire         rsp_xbar_demux_045_src0_endofpacket;                                                                // rsp_xbar_demux_045:src0_endofpacket -> rsp_xbar_mux_006:sink12_endofpacket
	wire         rsp_xbar_demux_045_src0_valid;                                                                      // rsp_xbar_demux_045:src0_valid -> rsp_xbar_mux_006:sink12_valid
	wire         rsp_xbar_demux_045_src0_startofpacket;                                                              // rsp_xbar_demux_045:src0_startofpacket -> rsp_xbar_mux_006:sink12_startofpacket
	wire  [94:0] rsp_xbar_demux_045_src0_data;                                                                       // rsp_xbar_demux_045:src0_data -> rsp_xbar_mux_006:sink12_data
	wire  [65:0] rsp_xbar_demux_045_src0_channel;                                                                    // rsp_xbar_demux_045:src0_channel -> rsp_xbar_mux_006:sink12_channel
	wire         rsp_xbar_demux_045_src0_ready;                                                                      // rsp_xbar_mux_006:sink12_ready -> rsp_xbar_demux_045:src0_ready
	wire         rsp_xbar_demux_046_src0_endofpacket;                                                                // rsp_xbar_demux_046:src0_endofpacket -> rsp_xbar_mux_006:sink13_endofpacket
	wire         rsp_xbar_demux_046_src0_valid;                                                                      // rsp_xbar_demux_046:src0_valid -> rsp_xbar_mux_006:sink13_valid
	wire         rsp_xbar_demux_046_src0_startofpacket;                                                              // rsp_xbar_demux_046:src0_startofpacket -> rsp_xbar_mux_006:sink13_startofpacket
	wire  [94:0] rsp_xbar_demux_046_src0_data;                                                                       // rsp_xbar_demux_046:src0_data -> rsp_xbar_mux_006:sink13_data
	wire  [65:0] rsp_xbar_demux_046_src0_channel;                                                                    // rsp_xbar_demux_046:src0_channel -> rsp_xbar_mux_006:sink13_channel
	wire         rsp_xbar_demux_046_src0_ready;                                                                      // rsp_xbar_mux_006:sink13_ready -> rsp_xbar_demux_046:src0_ready
	wire         rsp_xbar_demux_047_src0_endofpacket;                                                                // rsp_xbar_demux_047:src0_endofpacket -> rsp_xbar_mux_007:sink3_endofpacket
	wire         rsp_xbar_demux_047_src0_valid;                                                                      // rsp_xbar_demux_047:src0_valid -> rsp_xbar_mux_007:sink3_valid
	wire         rsp_xbar_demux_047_src0_startofpacket;                                                              // rsp_xbar_demux_047:src0_startofpacket -> rsp_xbar_mux_007:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_047_src0_data;                                                                       // rsp_xbar_demux_047:src0_data -> rsp_xbar_mux_007:sink3_data
	wire  [65:0] rsp_xbar_demux_047_src0_channel;                                                                    // rsp_xbar_demux_047:src0_channel -> rsp_xbar_mux_007:sink3_channel
	wire         rsp_xbar_demux_047_src0_ready;                                                                      // rsp_xbar_mux_007:sink3_ready -> rsp_xbar_demux_047:src0_ready
	wire         rsp_xbar_demux_048_src0_endofpacket;                                                                // rsp_xbar_demux_048:src0_endofpacket -> rsp_xbar_mux_007:sink4_endofpacket
	wire         rsp_xbar_demux_048_src0_valid;                                                                      // rsp_xbar_demux_048:src0_valid -> rsp_xbar_mux_007:sink4_valid
	wire         rsp_xbar_demux_048_src0_startofpacket;                                                              // rsp_xbar_demux_048:src0_startofpacket -> rsp_xbar_mux_007:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_048_src0_data;                                                                       // rsp_xbar_demux_048:src0_data -> rsp_xbar_mux_007:sink4_data
	wire  [65:0] rsp_xbar_demux_048_src0_channel;                                                                    // rsp_xbar_demux_048:src0_channel -> rsp_xbar_mux_007:sink4_channel
	wire         rsp_xbar_demux_048_src0_ready;                                                                      // rsp_xbar_mux_007:sink4_ready -> rsp_xbar_demux_048:src0_ready
	wire         rsp_xbar_demux_048_src1_endofpacket;                                                                // rsp_xbar_demux_048:src1_endofpacket -> rsp_xbar_mux_008:sink3_endofpacket
	wire         rsp_xbar_demux_048_src1_valid;                                                                      // rsp_xbar_demux_048:src1_valid -> rsp_xbar_mux_008:sink3_valid
	wire         rsp_xbar_demux_048_src1_startofpacket;                                                              // rsp_xbar_demux_048:src1_startofpacket -> rsp_xbar_mux_008:sink3_startofpacket
	wire  [94:0] rsp_xbar_demux_048_src1_data;                                                                       // rsp_xbar_demux_048:src1_data -> rsp_xbar_mux_008:sink3_data
	wire  [65:0] rsp_xbar_demux_048_src1_channel;                                                                    // rsp_xbar_demux_048:src1_channel -> rsp_xbar_mux_008:sink3_channel
	wire         rsp_xbar_demux_048_src1_ready;                                                                      // rsp_xbar_mux_008:sink3_ready -> rsp_xbar_demux_048:src1_ready
	wire         rsp_xbar_demux_049_src0_endofpacket;                                                                // rsp_xbar_demux_049:src0_endofpacket -> rsp_xbar_mux_007:sink5_endofpacket
	wire         rsp_xbar_demux_049_src0_valid;                                                                      // rsp_xbar_demux_049:src0_valid -> rsp_xbar_mux_007:sink5_valid
	wire         rsp_xbar_demux_049_src0_startofpacket;                                                              // rsp_xbar_demux_049:src0_startofpacket -> rsp_xbar_mux_007:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_049_src0_data;                                                                       // rsp_xbar_demux_049:src0_data -> rsp_xbar_mux_007:sink5_data
	wire  [65:0] rsp_xbar_demux_049_src0_channel;                                                                    // rsp_xbar_demux_049:src0_channel -> rsp_xbar_mux_007:sink5_channel
	wire         rsp_xbar_demux_049_src0_ready;                                                                      // rsp_xbar_mux_007:sink5_ready -> rsp_xbar_demux_049:src0_ready
	wire         rsp_xbar_demux_050_src0_endofpacket;                                                                // rsp_xbar_demux_050:src0_endofpacket -> rsp_xbar_mux_007:sink6_endofpacket
	wire         rsp_xbar_demux_050_src0_valid;                                                                      // rsp_xbar_demux_050:src0_valid -> rsp_xbar_mux_007:sink6_valid
	wire         rsp_xbar_demux_050_src0_startofpacket;                                                              // rsp_xbar_demux_050:src0_startofpacket -> rsp_xbar_mux_007:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_050_src0_data;                                                                       // rsp_xbar_demux_050:src0_data -> rsp_xbar_mux_007:sink6_data
	wire  [65:0] rsp_xbar_demux_050_src0_channel;                                                                    // rsp_xbar_demux_050:src0_channel -> rsp_xbar_mux_007:sink6_channel
	wire         rsp_xbar_demux_050_src0_ready;                                                                      // rsp_xbar_mux_007:sink6_ready -> rsp_xbar_demux_050:src0_ready
	wire         rsp_xbar_demux_051_src0_endofpacket;                                                                // rsp_xbar_demux_051:src0_endofpacket -> rsp_xbar_mux_007:sink7_endofpacket
	wire         rsp_xbar_demux_051_src0_valid;                                                                      // rsp_xbar_demux_051:src0_valid -> rsp_xbar_mux_007:sink7_valid
	wire         rsp_xbar_demux_051_src0_startofpacket;                                                              // rsp_xbar_demux_051:src0_startofpacket -> rsp_xbar_mux_007:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_051_src0_data;                                                                       // rsp_xbar_demux_051:src0_data -> rsp_xbar_mux_007:sink7_data
	wire  [65:0] rsp_xbar_demux_051_src0_channel;                                                                    // rsp_xbar_demux_051:src0_channel -> rsp_xbar_mux_007:sink7_channel
	wire         rsp_xbar_demux_051_src0_ready;                                                                      // rsp_xbar_mux_007:sink7_ready -> rsp_xbar_demux_051:src0_ready
	wire         rsp_xbar_demux_052_src0_endofpacket;                                                                // rsp_xbar_demux_052:src0_endofpacket -> rsp_xbar_mux_007:sink8_endofpacket
	wire         rsp_xbar_demux_052_src0_valid;                                                                      // rsp_xbar_demux_052:src0_valid -> rsp_xbar_mux_007:sink8_valid
	wire         rsp_xbar_demux_052_src0_startofpacket;                                                              // rsp_xbar_demux_052:src0_startofpacket -> rsp_xbar_mux_007:sink8_startofpacket
	wire  [94:0] rsp_xbar_demux_052_src0_data;                                                                       // rsp_xbar_demux_052:src0_data -> rsp_xbar_mux_007:sink8_data
	wire  [65:0] rsp_xbar_demux_052_src0_channel;                                                                    // rsp_xbar_demux_052:src0_channel -> rsp_xbar_mux_007:sink8_channel
	wire         rsp_xbar_demux_052_src0_ready;                                                                      // rsp_xbar_mux_007:sink8_ready -> rsp_xbar_demux_052:src0_ready
	wire         rsp_xbar_demux_052_src1_endofpacket;                                                                // rsp_xbar_demux_052:src1_endofpacket -> rsp_xbar_mux_008:sink4_endofpacket
	wire         rsp_xbar_demux_052_src1_valid;                                                                      // rsp_xbar_demux_052:src1_valid -> rsp_xbar_mux_008:sink4_valid
	wire         rsp_xbar_demux_052_src1_startofpacket;                                                              // rsp_xbar_demux_052:src1_startofpacket -> rsp_xbar_mux_008:sink4_startofpacket
	wire  [94:0] rsp_xbar_demux_052_src1_data;                                                                       // rsp_xbar_demux_052:src1_data -> rsp_xbar_mux_008:sink4_data
	wire  [65:0] rsp_xbar_demux_052_src1_channel;                                                                    // rsp_xbar_demux_052:src1_channel -> rsp_xbar_mux_008:sink4_channel
	wire         rsp_xbar_demux_052_src1_ready;                                                                      // rsp_xbar_mux_008:sink4_ready -> rsp_xbar_demux_052:src1_ready
	wire         rsp_xbar_demux_052_src2_endofpacket;                                                                // rsp_xbar_demux_052:src2_endofpacket -> rsp_xbar_mux_009:sink9_endofpacket
	wire         rsp_xbar_demux_052_src2_valid;                                                                      // rsp_xbar_demux_052:src2_valid -> rsp_xbar_mux_009:sink9_valid
	wire         rsp_xbar_demux_052_src2_startofpacket;                                                              // rsp_xbar_demux_052:src2_startofpacket -> rsp_xbar_mux_009:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_052_src2_data;                                                                       // rsp_xbar_demux_052:src2_data -> rsp_xbar_mux_009:sink9_data
	wire  [65:0] rsp_xbar_demux_052_src2_channel;                                                                    // rsp_xbar_demux_052:src2_channel -> rsp_xbar_mux_009:sink9_channel
	wire         rsp_xbar_demux_052_src2_ready;                                                                      // rsp_xbar_mux_009:sink9_ready -> rsp_xbar_demux_052:src2_ready
	wire         rsp_xbar_demux_052_src3_endofpacket;                                                                // rsp_xbar_demux_052:src3_endofpacket -> rsp_xbar_mux_010:sink9_endofpacket
	wire         rsp_xbar_demux_052_src3_valid;                                                                      // rsp_xbar_demux_052:src3_valid -> rsp_xbar_mux_010:sink9_valid
	wire         rsp_xbar_demux_052_src3_startofpacket;                                                              // rsp_xbar_demux_052:src3_startofpacket -> rsp_xbar_mux_010:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_052_src3_data;                                                                       // rsp_xbar_demux_052:src3_data -> rsp_xbar_mux_010:sink9_data
	wire  [65:0] rsp_xbar_demux_052_src3_channel;                                                                    // rsp_xbar_demux_052:src3_channel -> rsp_xbar_mux_010:sink9_channel
	wire         rsp_xbar_demux_052_src3_ready;                                                                      // rsp_xbar_mux_010:sink9_ready -> rsp_xbar_demux_052:src3_ready
	wire         rsp_xbar_demux_053_src0_endofpacket;                                                                // rsp_xbar_demux_053:src0_endofpacket -> rsp_xbar_mux_007:sink9_endofpacket
	wire         rsp_xbar_demux_053_src0_valid;                                                                      // rsp_xbar_demux_053:src0_valid -> rsp_xbar_mux_007:sink9_valid
	wire         rsp_xbar_demux_053_src0_startofpacket;                                                              // rsp_xbar_demux_053:src0_startofpacket -> rsp_xbar_mux_007:sink9_startofpacket
	wire  [94:0] rsp_xbar_demux_053_src0_data;                                                                       // rsp_xbar_demux_053:src0_data -> rsp_xbar_mux_007:sink9_data
	wire  [65:0] rsp_xbar_demux_053_src0_channel;                                                                    // rsp_xbar_demux_053:src0_channel -> rsp_xbar_mux_007:sink9_channel
	wire         rsp_xbar_demux_053_src0_ready;                                                                      // rsp_xbar_mux_007:sink9_ready -> rsp_xbar_demux_053:src0_ready
	wire         rsp_xbar_demux_053_src1_endofpacket;                                                                // rsp_xbar_demux_053:src1_endofpacket -> rsp_xbar_mux_008:sink5_endofpacket
	wire         rsp_xbar_demux_053_src1_valid;                                                                      // rsp_xbar_demux_053:src1_valid -> rsp_xbar_mux_008:sink5_valid
	wire         rsp_xbar_demux_053_src1_startofpacket;                                                              // rsp_xbar_demux_053:src1_startofpacket -> rsp_xbar_mux_008:sink5_startofpacket
	wire  [94:0] rsp_xbar_demux_053_src1_data;                                                                       // rsp_xbar_demux_053:src1_data -> rsp_xbar_mux_008:sink5_data
	wire  [65:0] rsp_xbar_demux_053_src1_channel;                                                                    // rsp_xbar_demux_053:src1_channel -> rsp_xbar_mux_008:sink5_channel
	wire         rsp_xbar_demux_053_src1_ready;                                                                      // rsp_xbar_mux_008:sink5_ready -> rsp_xbar_demux_053:src1_ready
	wire         rsp_xbar_demux_053_src2_endofpacket;                                                                // rsp_xbar_demux_053:src2_endofpacket -> rsp_xbar_mux_009:sink10_endofpacket
	wire         rsp_xbar_demux_053_src2_valid;                                                                      // rsp_xbar_demux_053:src2_valid -> rsp_xbar_mux_009:sink10_valid
	wire         rsp_xbar_demux_053_src2_startofpacket;                                                              // rsp_xbar_demux_053:src2_startofpacket -> rsp_xbar_mux_009:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_053_src2_data;                                                                       // rsp_xbar_demux_053:src2_data -> rsp_xbar_mux_009:sink10_data
	wire  [65:0] rsp_xbar_demux_053_src2_channel;                                                                    // rsp_xbar_demux_053:src2_channel -> rsp_xbar_mux_009:sink10_channel
	wire         rsp_xbar_demux_053_src2_ready;                                                                      // rsp_xbar_mux_009:sink10_ready -> rsp_xbar_demux_053:src2_ready
	wire         rsp_xbar_demux_053_src3_endofpacket;                                                                // rsp_xbar_demux_053:src3_endofpacket -> rsp_xbar_mux_010:sink10_endofpacket
	wire         rsp_xbar_demux_053_src3_valid;                                                                      // rsp_xbar_demux_053:src3_valid -> rsp_xbar_mux_010:sink10_valid
	wire         rsp_xbar_demux_053_src3_startofpacket;                                                              // rsp_xbar_demux_053:src3_startofpacket -> rsp_xbar_mux_010:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_053_src3_data;                                                                       // rsp_xbar_demux_053:src3_data -> rsp_xbar_mux_010:sink10_data
	wire  [65:0] rsp_xbar_demux_053_src3_channel;                                                                    // rsp_xbar_demux_053:src3_channel -> rsp_xbar_mux_010:sink10_channel
	wire         rsp_xbar_demux_053_src3_ready;                                                                      // rsp_xbar_mux_010:sink10_ready -> rsp_xbar_demux_053:src3_ready
	wire         rsp_xbar_demux_054_src0_endofpacket;                                                                // rsp_xbar_demux_054:src0_endofpacket -> rsp_xbar_mux_007:sink10_endofpacket
	wire         rsp_xbar_demux_054_src0_valid;                                                                      // rsp_xbar_demux_054:src0_valid -> rsp_xbar_mux_007:sink10_valid
	wire         rsp_xbar_demux_054_src0_startofpacket;                                                              // rsp_xbar_demux_054:src0_startofpacket -> rsp_xbar_mux_007:sink10_startofpacket
	wire  [94:0] rsp_xbar_demux_054_src0_data;                                                                       // rsp_xbar_demux_054:src0_data -> rsp_xbar_mux_007:sink10_data
	wire  [65:0] rsp_xbar_demux_054_src0_channel;                                                                    // rsp_xbar_demux_054:src0_channel -> rsp_xbar_mux_007:sink10_channel
	wire         rsp_xbar_demux_054_src0_ready;                                                                      // rsp_xbar_mux_007:sink10_ready -> rsp_xbar_demux_054:src0_ready
	wire         rsp_xbar_demux_054_src1_endofpacket;                                                                // rsp_xbar_demux_054:src1_endofpacket -> rsp_xbar_mux_008:sink6_endofpacket
	wire         rsp_xbar_demux_054_src1_valid;                                                                      // rsp_xbar_demux_054:src1_valid -> rsp_xbar_mux_008:sink6_valid
	wire         rsp_xbar_demux_054_src1_startofpacket;                                                              // rsp_xbar_demux_054:src1_startofpacket -> rsp_xbar_mux_008:sink6_startofpacket
	wire  [94:0] rsp_xbar_demux_054_src1_data;                                                                       // rsp_xbar_demux_054:src1_data -> rsp_xbar_mux_008:sink6_data
	wire  [65:0] rsp_xbar_demux_054_src1_channel;                                                                    // rsp_xbar_demux_054:src1_channel -> rsp_xbar_mux_008:sink6_channel
	wire         rsp_xbar_demux_054_src1_ready;                                                                      // rsp_xbar_mux_008:sink6_ready -> rsp_xbar_demux_054:src1_ready
	wire         rsp_xbar_demux_054_src2_endofpacket;                                                                // rsp_xbar_demux_054:src2_endofpacket -> rsp_xbar_mux_009:sink11_endofpacket
	wire         rsp_xbar_demux_054_src2_valid;                                                                      // rsp_xbar_demux_054:src2_valid -> rsp_xbar_mux_009:sink11_valid
	wire         rsp_xbar_demux_054_src2_startofpacket;                                                              // rsp_xbar_demux_054:src2_startofpacket -> rsp_xbar_mux_009:sink11_startofpacket
	wire  [94:0] rsp_xbar_demux_054_src2_data;                                                                       // rsp_xbar_demux_054:src2_data -> rsp_xbar_mux_009:sink11_data
	wire  [65:0] rsp_xbar_demux_054_src2_channel;                                                                    // rsp_xbar_demux_054:src2_channel -> rsp_xbar_mux_009:sink11_channel
	wire         rsp_xbar_demux_054_src2_ready;                                                                      // rsp_xbar_mux_009:sink11_ready -> rsp_xbar_demux_054:src2_ready
	wire         rsp_xbar_demux_054_src3_endofpacket;                                                                // rsp_xbar_demux_054:src3_endofpacket -> rsp_xbar_mux_010:sink11_endofpacket
	wire         rsp_xbar_demux_054_src3_valid;                                                                      // rsp_xbar_demux_054:src3_valid -> rsp_xbar_mux_010:sink11_valid
	wire         rsp_xbar_demux_054_src3_startofpacket;                                                              // rsp_xbar_demux_054:src3_startofpacket -> rsp_xbar_mux_010:sink11_startofpacket
	wire  [94:0] rsp_xbar_demux_054_src3_data;                                                                       // rsp_xbar_demux_054:src3_data -> rsp_xbar_mux_010:sink11_data
	wire  [65:0] rsp_xbar_demux_054_src3_channel;                                                                    // rsp_xbar_demux_054:src3_channel -> rsp_xbar_mux_010:sink11_channel
	wire         rsp_xbar_demux_054_src3_ready;                                                                      // rsp_xbar_mux_010:sink11_ready -> rsp_xbar_demux_054:src3_ready
	wire         rsp_xbar_demux_055_src0_endofpacket;                                                                // rsp_xbar_demux_055:src0_endofpacket -> rsp_xbar_mux_008:sink7_endofpacket
	wire         rsp_xbar_demux_055_src0_valid;                                                                      // rsp_xbar_demux_055:src0_valid -> rsp_xbar_mux_008:sink7_valid
	wire         rsp_xbar_demux_055_src0_startofpacket;                                                              // rsp_xbar_demux_055:src0_startofpacket -> rsp_xbar_mux_008:sink7_startofpacket
	wire  [94:0] rsp_xbar_demux_055_src0_data;                                                                       // rsp_xbar_demux_055:src0_data -> rsp_xbar_mux_008:sink7_data
	wire  [65:0] rsp_xbar_demux_055_src0_channel;                                                                    // rsp_xbar_demux_055:src0_channel -> rsp_xbar_mux_008:sink7_channel
	wire         rsp_xbar_demux_055_src0_ready;                                                                      // rsp_xbar_mux_008:sink7_ready -> rsp_xbar_demux_055:src0_ready
	wire         rsp_xbar_demux_056_src0_endofpacket;                                                                // rsp_xbar_demux_056:src0_endofpacket -> rsp_xbar_mux_009:sink12_endofpacket
	wire         rsp_xbar_demux_056_src0_valid;                                                                      // rsp_xbar_demux_056:src0_valid -> rsp_xbar_mux_009:sink12_valid
	wire         rsp_xbar_demux_056_src0_startofpacket;                                                              // rsp_xbar_demux_056:src0_startofpacket -> rsp_xbar_mux_009:sink12_startofpacket
	wire  [94:0] rsp_xbar_demux_056_src0_data;                                                                       // rsp_xbar_demux_056:src0_data -> rsp_xbar_mux_009:sink12_data
	wire  [65:0] rsp_xbar_demux_056_src0_channel;                                                                    // rsp_xbar_demux_056:src0_channel -> rsp_xbar_mux_009:sink12_channel
	wire         rsp_xbar_demux_056_src0_ready;                                                                      // rsp_xbar_mux_009:sink12_ready -> rsp_xbar_demux_056:src0_ready
	wire         rsp_xbar_demux_057_src0_endofpacket;                                                                // rsp_xbar_demux_057:src0_endofpacket -> rsp_xbar_mux_009:sink13_endofpacket
	wire         rsp_xbar_demux_057_src0_valid;                                                                      // rsp_xbar_demux_057:src0_valid -> rsp_xbar_mux_009:sink13_valid
	wire         rsp_xbar_demux_057_src0_startofpacket;                                                              // rsp_xbar_demux_057:src0_startofpacket -> rsp_xbar_mux_009:sink13_startofpacket
	wire  [94:0] rsp_xbar_demux_057_src0_data;                                                                       // rsp_xbar_demux_057:src0_data -> rsp_xbar_mux_009:sink13_data
	wire  [65:0] rsp_xbar_demux_057_src0_channel;                                                                    // rsp_xbar_demux_057:src0_channel -> rsp_xbar_mux_009:sink13_channel
	wire         rsp_xbar_demux_057_src0_ready;                                                                      // rsp_xbar_mux_009:sink13_ready -> rsp_xbar_demux_057:src0_ready
	wire         rsp_xbar_demux_057_src1_endofpacket;                                                                // rsp_xbar_demux_057:src1_endofpacket -> rsp_xbar_mux_010:sink12_endofpacket
	wire         rsp_xbar_demux_057_src1_valid;                                                                      // rsp_xbar_demux_057:src1_valid -> rsp_xbar_mux_010:sink12_valid
	wire         rsp_xbar_demux_057_src1_startofpacket;                                                              // rsp_xbar_demux_057:src1_startofpacket -> rsp_xbar_mux_010:sink12_startofpacket
	wire  [94:0] rsp_xbar_demux_057_src1_data;                                                                       // rsp_xbar_demux_057:src1_data -> rsp_xbar_mux_010:sink12_data
	wire  [65:0] rsp_xbar_demux_057_src1_channel;                                                                    // rsp_xbar_demux_057:src1_channel -> rsp_xbar_mux_010:sink12_channel
	wire         rsp_xbar_demux_057_src1_ready;                                                                      // rsp_xbar_mux_010:sink12_ready -> rsp_xbar_demux_057:src1_ready
	wire         rsp_xbar_demux_058_src0_endofpacket;                                                                // rsp_xbar_demux_058:src0_endofpacket -> rsp_xbar_mux_010:sink13_endofpacket
	wire         rsp_xbar_demux_058_src0_valid;                                                                      // rsp_xbar_demux_058:src0_valid -> rsp_xbar_mux_010:sink13_valid
	wire         rsp_xbar_demux_058_src0_startofpacket;                                                              // rsp_xbar_demux_058:src0_startofpacket -> rsp_xbar_mux_010:sink13_startofpacket
	wire  [94:0] rsp_xbar_demux_058_src0_data;                                                                       // rsp_xbar_demux_058:src0_data -> rsp_xbar_mux_010:sink13_data
	wire  [65:0] rsp_xbar_demux_058_src0_channel;                                                                    // rsp_xbar_demux_058:src0_channel -> rsp_xbar_mux_010:sink13_channel
	wire         rsp_xbar_demux_058_src0_ready;                                                                      // rsp_xbar_mux_010:sink13_ready -> rsp_xbar_demux_058:src0_ready
	wire         rsp_xbar_demux_059_src0_endofpacket;                                                                // rsp_xbar_demux_059:src0_endofpacket -> rsp_xbar_mux_010:sink14_endofpacket
	wire         rsp_xbar_demux_059_src0_valid;                                                                      // rsp_xbar_demux_059:src0_valid -> rsp_xbar_mux_010:sink14_valid
	wire         rsp_xbar_demux_059_src0_startofpacket;                                                              // rsp_xbar_demux_059:src0_startofpacket -> rsp_xbar_mux_010:sink14_startofpacket
	wire  [94:0] rsp_xbar_demux_059_src0_data;                                                                       // rsp_xbar_demux_059:src0_data -> rsp_xbar_mux_010:sink14_data
	wire  [65:0] rsp_xbar_demux_059_src0_channel;                                                                    // rsp_xbar_demux_059:src0_channel -> rsp_xbar_mux_010:sink14_channel
	wire         rsp_xbar_demux_059_src0_ready;                                                                      // rsp_xbar_mux_010:sink14_ready -> rsp_xbar_demux_059:src0_ready
	wire         rsp_xbar_demux_060_src0_endofpacket;                                                                // rsp_xbar_demux_060:src0_endofpacket -> rsp_xbar_mux_010:sink15_endofpacket
	wire         rsp_xbar_demux_060_src0_valid;                                                                      // rsp_xbar_demux_060:src0_valid -> rsp_xbar_mux_010:sink15_valid
	wire         rsp_xbar_demux_060_src0_startofpacket;                                                              // rsp_xbar_demux_060:src0_startofpacket -> rsp_xbar_mux_010:sink15_startofpacket
	wire  [94:0] rsp_xbar_demux_060_src0_data;                                                                       // rsp_xbar_demux_060:src0_data -> rsp_xbar_mux_010:sink15_data
	wire  [65:0] rsp_xbar_demux_060_src0_channel;                                                                    // rsp_xbar_demux_060:src0_channel -> rsp_xbar_mux_010:sink15_channel
	wire         rsp_xbar_demux_060_src0_ready;                                                                      // rsp_xbar_mux_010:sink15_ready -> rsp_xbar_demux_060:src0_ready
	wire         rsp_xbar_demux_061_src0_endofpacket;                                                                // rsp_xbar_demux_061:src0_endofpacket -> rsp_xbar_mux_010:sink16_endofpacket
	wire         rsp_xbar_demux_061_src0_valid;                                                                      // rsp_xbar_demux_061:src0_valid -> rsp_xbar_mux_010:sink16_valid
	wire         rsp_xbar_demux_061_src0_startofpacket;                                                              // rsp_xbar_demux_061:src0_startofpacket -> rsp_xbar_mux_010:sink16_startofpacket
	wire  [94:0] rsp_xbar_demux_061_src0_data;                                                                       // rsp_xbar_demux_061:src0_data -> rsp_xbar_mux_010:sink16_data
	wire  [65:0] rsp_xbar_demux_061_src0_channel;                                                                    // rsp_xbar_demux_061:src0_channel -> rsp_xbar_mux_010:sink16_channel
	wire         rsp_xbar_demux_061_src0_ready;                                                                      // rsp_xbar_mux_010:sink16_ready -> rsp_xbar_demux_061:src0_ready
	wire         rsp_xbar_demux_062_src0_endofpacket;                                                                // rsp_xbar_demux_062:src0_endofpacket -> rsp_xbar_mux_011:sink19_endofpacket
	wire         rsp_xbar_demux_062_src0_valid;                                                                      // rsp_xbar_demux_062:src0_valid -> rsp_xbar_mux_011:sink19_valid
	wire         rsp_xbar_demux_062_src0_startofpacket;                                                              // rsp_xbar_demux_062:src0_startofpacket -> rsp_xbar_mux_011:sink19_startofpacket
	wire  [94:0] rsp_xbar_demux_062_src0_data;                                                                       // rsp_xbar_demux_062:src0_data -> rsp_xbar_mux_011:sink19_data
	wire  [65:0] rsp_xbar_demux_062_src0_channel;                                                                    // rsp_xbar_demux_062:src0_channel -> rsp_xbar_mux_011:sink19_channel
	wire         rsp_xbar_demux_062_src0_ready;                                                                      // rsp_xbar_mux_011:sink19_ready -> rsp_xbar_demux_062:src0_ready
	wire         rsp_xbar_demux_063_src0_endofpacket;                                                                // rsp_xbar_demux_063:src0_endofpacket -> rsp_xbar_mux_011:sink20_endofpacket
	wire         rsp_xbar_demux_063_src0_valid;                                                                      // rsp_xbar_demux_063:src0_valid -> rsp_xbar_mux_011:sink20_valid
	wire         rsp_xbar_demux_063_src0_startofpacket;                                                              // rsp_xbar_demux_063:src0_startofpacket -> rsp_xbar_mux_011:sink20_startofpacket
	wire  [94:0] rsp_xbar_demux_063_src0_data;                                                                       // rsp_xbar_demux_063:src0_data -> rsp_xbar_mux_011:sink20_data
	wire  [65:0] rsp_xbar_demux_063_src0_channel;                                                                    // rsp_xbar_demux_063:src0_channel -> rsp_xbar_mux_011:sink20_channel
	wire         rsp_xbar_demux_063_src0_ready;                                                                      // rsp_xbar_mux_011:sink20_ready -> rsp_xbar_demux_063:src0_ready
	wire         rsp_xbar_demux_064_src0_endofpacket;                                                                // rsp_xbar_demux_064:src0_endofpacket -> rsp_xbar_mux_011:sink21_endofpacket
	wire         rsp_xbar_demux_064_src0_valid;                                                                      // rsp_xbar_demux_064:src0_valid -> rsp_xbar_mux_011:sink21_valid
	wire         rsp_xbar_demux_064_src0_startofpacket;                                                              // rsp_xbar_demux_064:src0_startofpacket -> rsp_xbar_mux_011:sink21_startofpacket
	wire  [94:0] rsp_xbar_demux_064_src0_data;                                                                       // rsp_xbar_demux_064:src0_data -> rsp_xbar_mux_011:sink21_data
	wire  [65:0] rsp_xbar_demux_064_src0_channel;                                                                    // rsp_xbar_demux_064:src0_channel -> rsp_xbar_mux_011:sink21_channel
	wire         rsp_xbar_demux_064_src0_ready;                                                                      // rsp_xbar_mux_011:sink21_ready -> rsp_xbar_demux_064:src0_ready
	wire         rsp_xbar_demux_065_src0_endofpacket;                                                                // rsp_xbar_demux_065:src0_endofpacket -> rsp_xbar_mux_011:sink22_endofpacket
	wire         rsp_xbar_demux_065_src0_valid;                                                                      // rsp_xbar_demux_065:src0_valid -> rsp_xbar_mux_011:sink22_valid
	wire         rsp_xbar_demux_065_src0_startofpacket;                                                              // rsp_xbar_demux_065:src0_startofpacket -> rsp_xbar_mux_011:sink22_startofpacket
	wire  [94:0] rsp_xbar_demux_065_src0_data;                                                                       // rsp_xbar_demux_065:src0_data -> rsp_xbar_mux_011:sink22_data
	wire  [65:0] rsp_xbar_demux_065_src0_channel;                                                                    // rsp_xbar_demux_065:src0_channel -> rsp_xbar_mux_011:sink22_channel
	wire         rsp_xbar_demux_065_src0_ready;                                                                      // rsp_xbar_mux_011:sink22_ready -> rsp_xbar_demux_065:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                        // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                      // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [94:0] limiter_cmd_src_data;                                                                               // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [65:0] limiter_cmd_src_channel;                                                                            // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                              // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                       // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                             // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                     // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [94:0] rsp_xbar_mux_src_data;                                                                              // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [65:0] rsp_xbar_mux_src_channel;                                                                           // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                             // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                    // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                  // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [94:0] limiter_001_cmd_src_data;                                                                           // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire  [65:0] limiter_001_cmd_src_channel;                                                                        // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                          // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                   // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                         // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                 // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [94:0] rsp_xbar_mux_001_src_data;                                                                          // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire  [65:0] rsp_xbar_mux_001_src_channel;                                                                       // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                         // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         addr_router_002_src_endofpacket;                                                                    // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire         addr_router_002_src_valid;                                                                          // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire         addr_router_002_src_startofpacket;                                                                  // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [94:0] addr_router_002_src_data;                                                                           // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire  [65:0] addr_router_002_src_channel;                                                                        // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire         addr_router_002_src_ready;                                                                          // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire         rsp_xbar_mux_002_src_endofpacket;                                                                   // rsp_xbar_mux_002:src_endofpacket -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_002_src_valid;                                                                         // rsp_xbar_mux_002:src_valid -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_002_src_startofpacket;                                                                 // rsp_xbar_mux_002:src_startofpacket -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] rsp_xbar_mux_002_src_data;                                                                          // rsp_xbar_mux_002:src_data -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] rsp_xbar_mux_002_src_channel;                                                                       // rsp_xbar_mux_002:src_channel -> cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_002_src_ready;                                                                         // cpu_5_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	wire         limiter_002_cmd_src_endofpacket;                                                                    // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire         limiter_002_cmd_src_startofpacket;                                                                  // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [94:0] limiter_002_cmd_src_data;                                                                           // limiter_002:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire  [65:0] limiter_002_cmd_src_channel;                                                                        // limiter_002:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire         limiter_002_cmd_src_ready;                                                                          // cmd_xbar_demux_003:sink_ready -> limiter_002:cmd_src_ready
	wire         rsp_xbar_mux_003_src_endofpacket;                                                                   // rsp_xbar_mux_003:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire         rsp_xbar_mux_003_src_valid;                                                                         // rsp_xbar_mux_003:src_valid -> limiter_002:rsp_sink_valid
	wire         rsp_xbar_mux_003_src_startofpacket;                                                                 // rsp_xbar_mux_003:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire  [94:0] rsp_xbar_mux_003_src_data;                                                                          // rsp_xbar_mux_003:src_data -> limiter_002:rsp_sink_data
	wire  [65:0] rsp_xbar_mux_003_src_channel;                                                                       // rsp_xbar_mux_003:src_channel -> limiter_002:rsp_sink_channel
	wire         rsp_xbar_mux_003_src_ready;                                                                         // limiter_002:rsp_sink_ready -> rsp_xbar_mux_003:src_ready
	wire         addr_router_004_src_endofpacket;                                                                    // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire         addr_router_004_src_valid;                                                                          // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire         addr_router_004_src_startofpacket;                                                                  // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [94:0] addr_router_004_src_data;                                                                           // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire  [65:0] addr_router_004_src_channel;                                                                        // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire         addr_router_004_src_ready;                                                                          // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire         rsp_xbar_mux_004_src_endofpacket;                                                                   // rsp_xbar_mux_004:src_endofpacket -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_004_src_valid;                                                                         // rsp_xbar_mux_004:src_valid -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_004_src_startofpacket;                                                                 // rsp_xbar_mux_004:src_startofpacket -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] rsp_xbar_mux_004_src_data;                                                                          // rsp_xbar_mux_004:src_data -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] rsp_xbar_mux_004_src_channel;                                                                       // rsp_xbar_mux_004:src_channel -> cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_004_src_ready;                                                                         // cpu_4_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_004:src_ready
	wire         limiter_003_cmd_src_endofpacket;                                                                    // limiter_003:cmd_src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire         limiter_003_cmd_src_startofpacket;                                                                  // limiter_003:cmd_src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [94:0] limiter_003_cmd_src_data;                                                                           // limiter_003:cmd_src_data -> cmd_xbar_demux_005:sink_data
	wire  [65:0] limiter_003_cmd_src_channel;                                                                        // limiter_003:cmd_src_channel -> cmd_xbar_demux_005:sink_channel
	wire         limiter_003_cmd_src_ready;                                                                          // cmd_xbar_demux_005:sink_ready -> limiter_003:cmd_src_ready
	wire         rsp_xbar_mux_005_src_endofpacket;                                                                   // rsp_xbar_mux_005:src_endofpacket -> limiter_003:rsp_sink_endofpacket
	wire         rsp_xbar_mux_005_src_valid;                                                                         // rsp_xbar_mux_005:src_valid -> limiter_003:rsp_sink_valid
	wire         rsp_xbar_mux_005_src_startofpacket;                                                                 // rsp_xbar_mux_005:src_startofpacket -> limiter_003:rsp_sink_startofpacket
	wire  [94:0] rsp_xbar_mux_005_src_data;                                                                          // rsp_xbar_mux_005:src_data -> limiter_003:rsp_sink_data
	wire  [65:0] rsp_xbar_mux_005_src_channel;                                                                       // rsp_xbar_mux_005:src_channel -> limiter_003:rsp_sink_channel
	wire         rsp_xbar_mux_005_src_ready;                                                                         // limiter_003:rsp_sink_ready -> rsp_xbar_mux_005:src_ready
	wire         addr_router_006_src_endofpacket;                                                                    // addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire         addr_router_006_src_valid;                                                                          // addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	wire         addr_router_006_src_startofpacket;                                                                  // addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire  [94:0] addr_router_006_src_data;                                                                           // addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	wire  [65:0] addr_router_006_src_channel;                                                                        // addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	wire         addr_router_006_src_ready;                                                                          // cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	wire         rsp_xbar_mux_006_src_endofpacket;                                                                   // rsp_xbar_mux_006:src_endofpacket -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_006_src_valid;                                                                         // rsp_xbar_mux_006:src_valid -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_006_src_startofpacket;                                                                 // rsp_xbar_mux_006:src_startofpacket -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] rsp_xbar_mux_006_src_data;                                                                          // rsp_xbar_mux_006:src_data -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] rsp_xbar_mux_006_src_channel;                                                                       // rsp_xbar_mux_006:src_channel -> cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_006_src_ready;                                                                         // cpu_3_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_006:src_ready
	wire         addr_router_007_src_endofpacket;                                                                    // addr_router_007:src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	wire         addr_router_007_src_valid;                                                                          // addr_router_007:src_valid -> cmd_xbar_demux_007:sink_valid
	wire         addr_router_007_src_startofpacket;                                                                  // addr_router_007:src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	wire  [94:0] addr_router_007_src_data;                                                                           // addr_router_007:src_data -> cmd_xbar_demux_007:sink_data
	wire  [65:0] addr_router_007_src_channel;                                                                        // addr_router_007:src_channel -> cmd_xbar_demux_007:sink_channel
	wire         addr_router_007_src_ready;                                                                          // cmd_xbar_demux_007:sink_ready -> addr_router_007:src_ready
	wire         rsp_xbar_mux_007_src_endofpacket;                                                                   // rsp_xbar_mux_007:src_endofpacket -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_007_src_valid;                                                                         // rsp_xbar_mux_007:src_valid -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_007_src_startofpacket;                                                                 // rsp_xbar_mux_007:src_startofpacket -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] rsp_xbar_mux_007_src_data;                                                                          // rsp_xbar_mux_007:src_data -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] rsp_xbar_mux_007_src_channel;                                                                       // rsp_xbar_mux_007:src_channel -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_007_src_ready;                                                                         // cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_007:src_ready
	wire         limiter_004_cmd_src_endofpacket;                                                                    // limiter_004:cmd_src_endofpacket -> cmd_xbar_demux_008:sink_endofpacket
	wire         limiter_004_cmd_src_startofpacket;                                                                  // limiter_004:cmd_src_startofpacket -> cmd_xbar_demux_008:sink_startofpacket
	wire  [94:0] limiter_004_cmd_src_data;                                                                           // limiter_004:cmd_src_data -> cmd_xbar_demux_008:sink_data
	wire  [65:0] limiter_004_cmd_src_channel;                                                                        // limiter_004:cmd_src_channel -> cmd_xbar_demux_008:sink_channel
	wire         limiter_004_cmd_src_ready;                                                                          // cmd_xbar_demux_008:sink_ready -> limiter_004:cmd_src_ready
	wire         rsp_xbar_mux_008_src_endofpacket;                                                                   // rsp_xbar_mux_008:src_endofpacket -> limiter_004:rsp_sink_endofpacket
	wire         rsp_xbar_mux_008_src_valid;                                                                         // rsp_xbar_mux_008:src_valid -> limiter_004:rsp_sink_valid
	wire         rsp_xbar_mux_008_src_startofpacket;                                                                 // rsp_xbar_mux_008:src_startofpacket -> limiter_004:rsp_sink_startofpacket
	wire  [94:0] rsp_xbar_mux_008_src_data;                                                                          // rsp_xbar_mux_008:src_data -> limiter_004:rsp_sink_data
	wire  [65:0] rsp_xbar_mux_008_src_channel;                                                                       // rsp_xbar_mux_008:src_channel -> limiter_004:rsp_sink_channel
	wire         rsp_xbar_mux_008_src_ready;                                                                         // limiter_004:rsp_sink_ready -> rsp_xbar_mux_008:src_ready
	wire         limiter_005_cmd_src_endofpacket;                                                                    // limiter_005:cmd_src_endofpacket -> cmd_xbar_demux_009:sink_endofpacket
	wire         limiter_005_cmd_src_startofpacket;                                                                  // limiter_005:cmd_src_startofpacket -> cmd_xbar_demux_009:sink_startofpacket
	wire  [94:0] limiter_005_cmd_src_data;                                                                           // limiter_005:cmd_src_data -> cmd_xbar_demux_009:sink_data
	wire  [65:0] limiter_005_cmd_src_channel;                                                                        // limiter_005:cmd_src_channel -> cmd_xbar_demux_009:sink_channel
	wire         limiter_005_cmd_src_ready;                                                                          // cmd_xbar_demux_009:sink_ready -> limiter_005:cmd_src_ready
	wire         rsp_xbar_mux_009_src_endofpacket;                                                                   // rsp_xbar_mux_009:src_endofpacket -> limiter_005:rsp_sink_endofpacket
	wire         rsp_xbar_mux_009_src_valid;                                                                         // rsp_xbar_mux_009:src_valid -> limiter_005:rsp_sink_valid
	wire         rsp_xbar_mux_009_src_startofpacket;                                                                 // rsp_xbar_mux_009:src_startofpacket -> limiter_005:rsp_sink_startofpacket
	wire  [94:0] rsp_xbar_mux_009_src_data;                                                                          // rsp_xbar_mux_009:src_data -> limiter_005:rsp_sink_data
	wire  [65:0] rsp_xbar_mux_009_src_channel;                                                                       // rsp_xbar_mux_009:src_channel -> limiter_005:rsp_sink_channel
	wire         rsp_xbar_mux_009_src_ready;                                                                         // limiter_005:rsp_sink_ready -> rsp_xbar_mux_009:src_ready
	wire         addr_router_010_src_endofpacket;                                                                    // addr_router_010:src_endofpacket -> cmd_xbar_demux_010:sink_endofpacket
	wire         addr_router_010_src_valid;                                                                          // addr_router_010:src_valid -> cmd_xbar_demux_010:sink_valid
	wire         addr_router_010_src_startofpacket;                                                                  // addr_router_010:src_startofpacket -> cmd_xbar_demux_010:sink_startofpacket
	wire  [94:0] addr_router_010_src_data;                                                                           // addr_router_010:src_data -> cmd_xbar_demux_010:sink_data
	wire  [65:0] addr_router_010_src_channel;                                                                        // addr_router_010:src_channel -> cmd_xbar_demux_010:sink_channel
	wire         addr_router_010_src_ready;                                                                          // cmd_xbar_demux_010:sink_ready -> addr_router_010:src_ready
	wire         rsp_xbar_mux_010_src_endofpacket;                                                                   // rsp_xbar_mux_010:src_endofpacket -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_010_src_valid;                                                                         // rsp_xbar_mux_010:src_valid -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_010_src_startofpacket;                                                                 // rsp_xbar_mux_010:src_startofpacket -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] rsp_xbar_mux_010_src_data;                                                                          // rsp_xbar_mux_010:src_data -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] rsp_xbar_mux_010_src_channel;                                                                       // rsp_xbar_mux_010:src_channel -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_010_src_ready;                                                                         // cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_010:src_ready
	wire         addr_router_011_src_endofpacket;                                                                    // addr_router_011:src_endofpacket -> cmd_xbar_demux_011:sink_endofpacket
	wire         addr_router_011_src_valid;                                                                          // addr_router_011:src_valid -> cmd_xbar_demux_011:sink_valid
	wire         addr_router_011_src_startofpacket;                                                                  // addr_router_011:src_startofpacket -> cmd_xbar_demux_011:sink_startofpacket
	wire  [94:0] addr_router_011_src_data;                                                                           // addr_router_011:src_data -> cmd_xbar_demux_011:sink_data
	wire  [65:0] addr_router_011_src_channel;                                                                        // addr_router_011:src_channel -> cmd_xbar_demux_011:sink_channel
	wire         addr_router_011_src_ready;                                                                          // cmd_xbar_demux_011:sink_ready -> addr_router_011:src_ready
	wire         rsp_xbar_mux_011_src_endofpacket;                                                                   // rsp_xbar_mux_011:src_endofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_011_src_valid;                                                                         // rsp_xbar_mux_011:src_valid -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_011_src_startofpacket;                                                                 // rsp_xbar_mux_011:src_startofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] rsp_xbar_mux_011_src_data;                                                                          // rsp_xbar_mux_011:src_data -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [65:0] rsp_xbar_mux_011_src_channel;                                                                       // rsp_xbar_mux_011:src_channel -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_011_src_ready;                                                                         // cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_011:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                       // cmd_xbar_mux:src_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                             // cmd_xbar_mux:src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                     // cmd_xbar_mux:src_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_src_data;                                                                              // cmd_xbar_mux:src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_src_channel;                                                                           // cmd_xbar_mux:src_channel -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                          // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                        // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [94:0] id_router_src_data;                                                                                 // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [65:0] id_router_src_channel;                                                                              // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                                          // ins_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                                      // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                            // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                    // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [94:0] id_router_001_src_data;                                                                             // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [65:0] id_router_001_src_channel;                                                                          // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                   // cmd_xbar_mux_002:src_endofpacket -> atob_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                         // cmd_xbar_mux_002:src_valid -> atob_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                 // cmd_xbar_mux_002:src_startofpacket -> atob_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_002_src_data;                                                                          // cmd_xbar_mux_002:src_data -> atob_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_002_src_channel;                                                                       // cmd_xbar_mux_002:src_channel -> atob_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                         // atob_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                      // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                            // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                    // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [94:0] id_router_002_src_data;                                                                             // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [65:0] id_router_002_src_channel;                                                                          // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                   // cmd_xbar_mux_003:src_endofpacket -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                         // cmd_xbar_mux_003:src_valid -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                                 // cmd_xbar_mux_003:src_startofpacket -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_003_src_data;                                                                          // cmd_xbar_mux_003:src_data -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_003_src_channel;                                                                       // cmd_xbar_mux_003:src_channel -> atob_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                         // atob_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire         id_router_003_src_endofpacket;                                                                      // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                            // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                    // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [94:0] id_router_003_src_data;                                                                             // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [65:0] id_router_003_src_channel;                                                                          // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_mux_004_src_endofpacket;                                                                   // cmd_xbar_mux_004:src_endofpacket -> atob_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_004_src_valid;                                                                         // cmd_xbar_mux_004:src_valid -> atob_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_004_src_startofpacket;                                                                 // cmd_xbar_mux_004:src_startofpacket -> atob_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_004_src_data;                                                                          // cmd_xbar_mux_004:src_data -> atob_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_004_src_channel;                                                                       // cmd_xbar_mux_004:src_channel -> atob_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_004_src_ready;                                                                         // atob_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire         id_router_004_src_endofpacket;                                                                      // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                            // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                    // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [94:0] id_router_004_src_data;                                                                             // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [65:0] id_router_004_src_channel;                                                                          // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_mux_005_src_endofpacket;                                                                   // cmd_xbar_mux_005:src_endofpacket -> atob_1_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_005_src_valid;                                                                         // cmd_xbar_mux_005:src_valid -> atob_1_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_005_src_startofpacket;                                                                 // cmd_xbar_mux_005:src_startofpacket -> atob_1_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_005_src_data;                                                                          // cmd_xbar_mux_005:src_data -> atob_1_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_005_src_channel;                                                                       // cmd_xbar_mux_005:src_channel -> atob_1_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_005_src_ready;                                                                         // atob_1_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire         id_router_005_src_endofpacket;                                                                      // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                            // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                    // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [94:0] id_router_005_src_data;                                                                             // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [65:0] id_router_005_src_channel;                                                                          // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                            // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_mux_006_src_endofpacket;                                                                   // cmd_xbar_mux_006:src_endofpacket -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_006_src_valid;                                                                         // cmd_xbar_mux_006:src_valid -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_006_src_startofpacket;                                                                 // cmd_xbar_mux_006:src_startofpacket -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_006_src_data;                                                                          // cmd_xbar_mux_006:src_data -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_006_src_channel;                                                                       // cmd_xbar_mux_006:src_channel -> atob_1_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_006_src_ready;                                                                         // atob_1_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	wire         id_router_006_src_endofpacket;                                                                      // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                            // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                    // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [94:0] id_router_006_src_data;                                                                             // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [65:0] id_router_006_src_channel;                                                                          // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                            // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_mux_007_src_endofpacket;                                                                   // cmd_xbar_mux_007:src_endofpacket -> atob_1_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_007_src_valid;                                                                         // cmd_xbar_mux_007:src_valid -> atob_1_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_007_src_startofpacket;                                                                 // cmd_xbar_mux_007:src_startofpacket -> atob_1_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_007_src_data;                                                                          // cmd_xbar_mux_007:src_data -> atob_1_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_007_src_channel;                                                                       // cmd_xbar_mux_007:src_channel -> atob_1_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_007_src_ready;                                                                         // atob_1_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	wire         id_router_007_src_endofpacket;                                                                      // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                            // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                    // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [94:0] id_router_007_src_data;                                                                             // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [65:0] id_router_007_src_channel;                                                                          // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                            // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_mux_008_src_endofpacket;                                                                   // cmd_xbar_mux_008:src_endofpacket -> atob_2_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_008_src_valid;                                                                         // cmd_xbar_mux_008:src_valid -> atob_2_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_008_src_startofpacket;                                                                 // cmd_xbar_mux_008:src_startofpacket -> atob_2_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_008_src_data;                                                                          // cmd_xbar_mux_008:src_data -> atob_2_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_008_src_channel;                                                                       // cmd_xbar_mux_008:src_channel -> atob_2_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_008_src_ready;                                                                         // atob_2_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire         id_router_008_src_endofpacket;                                                                      // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                            // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                    // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [94:0] id_router_008_src_data;                                                                             // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [65:0] id_router_008_src_channel;                                                                          // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                            // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_mux_009_src_endofpacket;                                                                   // cmd_xbar_mux_009:src_endofpacket -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_009_src_valid;                                                                         // cmd_xbar_mux_009:src_valid -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_009_src_startofpacket;                                                                 // cmd_xbar_mux_009:src_startofpacket -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_009_src_data;                                                                          // cmd_xbar_mux_009:src_data -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_009_src_channel;                                                                       // cmd_xbar_mux_009:src_channel -> atob_2_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_009_src_ready;                                                                         // atob_2_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire         id_router_009_src_endofpacket;                                                                      // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                            // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                    // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [94:0] id_router_009_src_data;                                                                             // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [65:0] id_router_009_src_channel;                                                                          // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                            // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_mux_010_src_endofpacket;                                                                   // cmd_xbar_mux_010:src_endofpacket -> atob_2_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_010_src_valid;                                                                         // cmd_xbar_mux_010:src_valid -> atob_2_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_010_src_startofpacket;                                                                 // cmd_xbar_mux_010:src_startofpacket -> atob_2_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_010_src_data;                                                                          // cmd_xbar_mux_010:src_data -> atob_2_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_010_src_channel;                                                                       // cmd_xbar_mux_010:src_channel -> atob_2_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_010_src_ready;                                                                         // atob_2_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire         id_router_010_src_endofpacket;                                                                      // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                            // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                    // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [94:0] id_router_010_src_data;                                                                             // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [65:0] id_router_010_src_channel;                                                                          // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                            // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_mux_011_src_endofpacket;                                                                   // cmd_xbar_mux_011:src_endofpacket -> atod_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_011_src_valid;                                                                         // cmd_xbar_mux_011:src_valid -> atod_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_011_src_startofpacket;                                                                 // cmd_xbar_mux_011:src_startofpacket -> atod_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_011_src_data;                                                                          // cmd_xbar_mux_011:src_data -> atod_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_011_src_channel;                                                                       // cmd_xbar_mux_011:src_channel -> atod_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_011_src_ready;                                                                         // atod_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_011:src_ready
	wire         id_router_011_src_endofpacket;                                                                      // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                            // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                    // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [94:0] id_router_011_src_data;                                                                             // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [65:0] id_router_011_src_channel;                                                                          // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                            // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_mux_012_src_endofpacket;                                                                   // cmd_xbar_mux_012:src_endofpacket -> atod_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_012_src_valid;                                                                         // cmd_xbar_mux_012:src_valid -> atod_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_012_src_startofpacket;                                                                 // cmd_xbar_mux_012:src_startofpacket -> atod_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_012_src_data;                                                                          // cmd_xbar_mux_012:src_data -> atod_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_012_src_channel;                                                                       // cmd_xbar_mux_012:src_channel -> atod_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_012_src_ready;                                                                         // atod_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_012:src_ready
	wire         id_router_012_src_endofpacket;                                                                      // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                            // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                    // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [94:0] id_router_012_src_data;                                                                             // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [65:0] id_router_012_src_channel;                                                                          // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                            // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_mux_013_src_endofpacket;                                                                   // cmd_xbar_mux_013:src_endofpacket -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_013_src_valid;                                                                         // cmd_xbar_mux_013:src_valid -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_013_src_startofpacket;                                                                 // cmd_xbar_mux_013:src_startofpacket -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_013_src_data;                                                                          // cmd_xbar_mux_013:src_data -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_013_src_channel;                                                                       // cmd_xbar_mux_013:src_channel -> atod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_013_src_ready;                                                                         // atod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	wire         id_router_013_src_endofpacket;                                                                      // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                            // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                    // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [94:0] id_router_013_src_data;                                                                             // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire  [65:0] id_router_013_src_channel;                                                                          // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                            // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire         cmd_xbar_mux_014_src_endofpacket;                                                                   // cmd_xbar_mux_014:src_endofpacket -> atoe_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_014_src_valid;                                                                         // cmd_xbar_mux_014:src_valid -> atoe_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_014_src_startofpacket;                                                                 // cmd_xbar_mux_014:src_startofpacket -> atoe_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_014_src_data;                                                                          // cmd_xbar_mux_014:src_data -> atoe_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_014_src_channel;                                                                       // cmd_xbar_mux_014:src_channel -> atoe_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_014_src_ready;                                                                         // atoe_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_014:src_ready
	wire         id_router_014_src_endofpacket;                                                                      // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire         id_router_014_src_valid;                                                                            // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire         id_router_014_src_startofpacket;                                                                    // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [94:0] id_router_014_src_data;                                                                             // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire  [65:0] id_router_014_src_channel;                                                                          // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire         id_router_014_src_ready;                                                                            // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire         cmd_xbar_mux_015_src_endofpacket;                                                                   // cmd_xbar_mux_015:src_endofpacket -> atoe_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_015_src_valid;                                                                         // cmd_xbar_mux_015:src_valid -> atoe_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_015_src_startofpacket;                                                                 // cmd_xbar_mux_015:src_startofpacket -> atoe_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_015_src_data;                                                                          // cmd_xbar_mux_015:src_data -> atoe_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_015_src_channel;                                                                       // cmd_xbar_mux_015:src_channel -> atoe_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_015_src_ready;                                                                         // atoe_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_015:src_ready
	wire         id_router_015_src_endofpacket;                                                                      // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire         id_router_015_src_valid;                                                                            // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire         id_router_015_src_startofpacket;                                                                    // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [94:0] id_router_015_src_data;                                                                             // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire  [65:0] id_router_015_src_channel;                                                                          // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire         id_router_015_src_ready;                                                                            // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire         cmd_xbar_mux_016_src_endofpacket;                                                                   // cmd_xbar_mux_016:src_endofpacket -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_016_src_valid;                                                                         // cmd_xbar_mux_016:src_valid -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_016_src_startofpacket;                                                                 // cmd_xbar_mux_016:src_startofpacket -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_016_src_data;                                                                          // cmd_xbar_mux_016:src_data -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_016_src_channel;                                                                       // cmd_xbar_mux_016:src_channel -> atoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_016_src_ready;                                                                         // atoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_016:src_ready
	wire         id_router_016_src_endofpacket;                                                                      // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire         id_router_016_src_valid;                                                                            // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire         id_router_016_src_startofpacket;                                                                    // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [94:0] id_router_016_src_data;                                                                             // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire  [65:0] id_router_016_src_channel;                                                                          // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire         id_router_016_src_ready;                                                                            // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire         cmd_xbar_mux_017_src_endofpacket;                                                                   // cmd_xbar_mux_017:src_endofpacket -> atof_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_017_src_valid;                                                                         // cmd_xbar_mux_017:src_valid -> atof_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_017_src_startofpacket;                                                                 // cmd_xbar_mux_017:src_startofpacket -> atof_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_017_src_data;                                                                          // cmd_xbar_mux_017:src_data -> atof_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_017_src_channel;                                                                       // cmd_xbar_mux_017:src_channel -> atof_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_017_src_ready;                                                                         // atof_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_017:src_ready
	wire         id_router_017_src_endofpacket;                                                                      // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire         id_router_017_src_valid;                                                                            // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire         id_router_017_src_startofpacket;                                                                    // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [94:0] id_router_017_src_data;                                                                             // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire  [65:0] id_router_017_src_channel;                                                                          // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire         id_router_017_src_ready;                                                                            // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire         cmd_xbar_mux_018_src_endofpacket;                                                                   // cmd_xbar_mux_018:src_endofpacket -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_018_src_valid;                                                                         // cmd_xbar_mux_018:src_valid -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_018_src_startofpacket;                                                                 // cmd_xbar_mux_018:src_startofpacket -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_018_src_data;                                                                          // cmd_xbar_mux_018:src_data -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_018_src_channel;                                                                       // cmd_xbar_mux_018:src_channel -> atof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_018_src_ready;                                                                         // atof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_018:src_ready
	wire         id_router_018_src_endofpacket;                                                                      // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire         id_router_018_src_valid;                                                                            // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire         id_router_018_src_startofpacket;                                                                    // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [94:0] id_router_018_src_data;                                                                             // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire  [65:0] id_router_018_src_channel;                                                                          // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire         id_router_018_src_ready;                                                                            // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire         cmd_xbar_mux_019_src_endofpacket;                                                                   // cmd_xbar_mux_019:src_endofpacket -> atof_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_019_src_valid;                                                                         // cmd_xbar_mux_019:src_valid -> atof_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_019_src_startofpacket;                                                                 // cmd_xbar_mux_019:src_startofpacket -> atof_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_019_src_data;                                                                          // cmd_xbar_mux_019:src_data -> atof_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_019_src_channel;                                                                       // cmd_xbar_mux_019:src_channel -> atof_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_019_src_ready;                                                                         // atof_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_019:src_ready
	wire         id_router_019_src_endofpacket;                                                                      // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire         id_router_019_src_valid;                                                                            // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire         id_router_019_src_startofpacket;                                                                    // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [94:0] id_router_019_src_data;                                                                             // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire  [65:0] id_router_019_src_channel;                                                                          // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire         id_router_019_src_ready;                                                                            // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                      // ins_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_020_src_endofpacket;                                                                      // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire         id_router_020_src_valid;                                                                            // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire         id_router_020_src_startofpacket;                                                                    // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [94:0] id_router_020_src_data;                                                                             // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire  [65:0] id_router_020_src_channel;                                                                          // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire         id_router_020_src_ready;                                                                            // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire         cmd_xbar_mux_021_src_endofpacket;                                                                   // cmd_xbar_mux_021:src_endofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_021_src_valid;                                                                         // cmd_xbar_mux_021:src_valid -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_021_src_startofpacket;                                                                 // cmd_xbar_mux_021:src_startofpacket -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_021_src_data;                                                                          // cmd_xbar_mux_021:src_data -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_021_src_channel;                                                                       // cmd_xbar_mux_021:src_channel -> cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_021_src_ready;                                                                         // cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_021:src_ready
	wire         id_router_021_src_endofpacket;                                                                      // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire         id_router_021_src_valid;                                                                            // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire         id_router_021_src_startofpacket;                                                                    // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [94:0] id_router_021_src_data;                                                                             // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire  [65:0] id_router_021_src_channel;                                                                          // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire         id_router_021_src_ready;                                                                            // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire         cmd_xbar_mux_022_src_endofpacket;                                                                   // cmd_xbar_mux_022:src_endofpacket -> etof_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_022_src_valid;                                                                         // cmd_xbar_mux_022:src_valid -> etof_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_022_src_startofpacket;                                                                 // cmd_xbar_mux_022:src_startofpacket -> etof_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_022_src_data;                                                                          // cmd_xbar_mux_022:src_data -> etof_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_022_src_channel;                                                                       // cmd_xbar_mux_022:src_channel -> etof_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_022_src_ready;                                                                         // etof_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_022:src_ready
	wire         id_router_022_src_endofpacket;                                                                      // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire         id_router_022_src_valid;                                                                            // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire         id_router_022_src_startofpacket;                                                                    // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [94:0] id_router_022_src_data;                                                                             // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire  [65:0] id_router_022_src_channel;                                                                          // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire         id_router_022_src_ready;                                                                            // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire         cmd_xbar_mux_023_src_endofpacket;                                                                   // cmd_xbar_mux_023:src_endofpacket -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_023_src_valid;                                                                         // cmd_xbar_mux_023:src_valid -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_023_src_startofpacket;                                                                 // cmd_xbar_mux_023:src_startofpacket -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_023_src_data;                                                                          // cmd_xbar_mux_023:src_data -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_023_src_channel;                                                                       // cmd_xbar_mux_023:src_channel -> etof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_023_src_ready;                                                                         // etof_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_023:src_ready
	wire         id_router_023_src_endofpacket;                                                                      // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire         id_router_023_src_valid;                                                                            // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire         id_router_023_src_startofpacket;                                                                    // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [94:0] id_router_023_src_data;                                                                             // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire  [65:0] id_router_023_src_channel;                                                                          // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire         id_router_023_src_ready;                                                                            // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire         cmd_xbar_mux_024_src_endofpacket;                                                                   // cmd_xbar_mux_024:src_endofpacket -> etof_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_024_src_valid;                                                                         // cmd_xbar_mux_024:src_valid -> etof_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_024_src_startofpacket;                                                                 // cmd_xbar_mux_024:src_startofpacket -> etof_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_024_src_data;                                                                          // cmd_xbar_mux_024:src_data -> etof_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_024_src_channel;                                                                       // cmd_xbar_mux_024:src_channel -> etof_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_024_src_ready;                                                                         // etof_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_024:src_ready
	wire         id_router_024_src_endofpacket;                                                                      // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire         id_router_024_src_valid;                                                                            // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire         id_router_024_src_startofpacket;                                                                    // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [94:0] id_router_024_src_data;                                                                             // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire  [65:0] id_router_024_src_channel;                                                                          // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire         id_router_024_src_ready;                                                                            // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire         cmd_xbar_demux_002_src7_ready;                                                                      // data_mem_5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src7_ready
	wire         id_router_025_src_endofpacket;                                                                      // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire         id_router_025_src_valid;                                                                            // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire         id_router_025_src_startofpacket;                                                                    // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire  [94:0] id_router_025_src_data;                                                                             // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire  [65:0] id_router_025_src_channel;                                                                          // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire         id_router_025_src_ready;                                                                            // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire         cmd_xbar_demux_002_src8_ready;                                                                      // jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src8_ready
	wire         id_router_026_src_endofpacket;                                                                      // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire         id_router_026_src_valid;                                                                            // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire         id_router_026_src_startofpacket;                                                                    // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire  [94:0] id_router_026_src_data;                                                                             // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire  [65:0] id_router_026_src_channel;                                                                          // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire         id_router_026_src_ready;                                                                            // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire         cmd_xbar_demux_002_src9_ready;                                                                      // timer_5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src9_ready
	wire         id_router_027_src_endofpacket;                                                                      // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire         id_router_027_src_valid;                                                                            // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire         id_router_027_src_startofpacket;                                                                    // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire  [94:0] id_router_027_src_data;                                                                             // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire  [65:0] id_router_027_src_channel;                                                                          // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire         id_router_027_src_ready;                                                                            // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire         cmd_xbar_demux_002_src10_ready;                                                                     // high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src10_ready
	wire         id_router_028_src_endofpacket;                                                                      // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire         id_router_028_src_valid;                                                                            // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire         id_router_028_src_startofpacket;                                                                    // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire  [94:0] id_router_028_src_data;                                                                             // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire  [65:0] id_router_028_src_channel;                                                                          // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire         id_router_028_src_ready;                                                                            // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire         cmd_xbar_demux_003_src6_ready;                                                                      // ins_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src6_ready
	wire         id_router_029_src_endofpacket;                                                                      // id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire         id_router_029_src_valid;                                                                            // id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	wire         id_router_029_src_startofpacket;                                                                    // id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire  [94:0] id_router_029_src_data;                                                                             // id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	wire  [65:0] id_router_029_src_channel;                                                                          // id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	wire         id_router_029_src_ready;                                                                            // rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	wire         cmd_xbar_mux_030_src_endofpacket;                                                                   // cmd_xbar_mux_030:src_endofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_030_src_valid;                                                                         // cmd_xbar_mux_030:src_valid -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_030_src_startofpacket;                                                                 // cmd_xbar_mux_030:src_startofpacket -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_030_src_data;                                                                          // cmd_xbar_mux_030:src_data -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_030_src_channel;                                                                       // cmd_xbar_mux_030:src_channel -> cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_030_src_ready;                                                                         // cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_030:src_ready
	wire         id_router_030_src_endofpacket;                                                                      // id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire         id_router_030_src_valid;                                                                            // id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	wire         id_router_030_src_startofpacket;                                                                    // id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire  [94:0] id_router_030_src_data;                                                                             // id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	wire  [65:0] id_router_030_src_channel;                                                                          // id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	wire         id_router_030_src_ready;                                                                            // rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	wire         cmd_xbar_mux_031_src_endofpacket;                                                                   // cmd_xbar_mux_031:src_endofpacket -> dtoe_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_031_src_valid;                                                                         // cmd_xbar_mux_031:src_valid -> dtoe_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_031_src_startofpacket;                                                                 // cmd_xbar_mux_031:src_startofpacket -> dtoe_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_031_src_data;                                                                          // cmd_xbar_mux_031:src_data -> dtoe_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_031_src_channel;                                                                       // cmd_xbar_mux_031:src_channel -> dtoe_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_031_src_ready;                                                                         // dtoe_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_031:src_ready
	wire         id_router_031_src_endofpacket;                                                                      // id_router_031:src_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	wire         id_router_031_src_valid;                                                                            // id_router_031:src_valid -> rsp_xbar_demux_031:sink_valid
	wire         id_router_031_src_startofpacket;                                                                    // id_router_031:src_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	wire  [94:0] id_router_031_src_data;                                                                             // id_router_031:src_data -> rsp_xbar_demux_031:sink_data
	wire  [65:0] id_router_031_src_channel;                                                                          // id_router_031:src_channel -> rsp_xbar_demux_031:sink_channel
	wire         id_router_031_src_ready;                                                                            // rsp_xbar_demux_031:sink_ready -> id_router_031:src_ready
	wire         cmd_xbar_mux_032_src_endofpacket;                                                                   // cmd_xbar_mux_032:src_endofpacket -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_032_src_valid;                                                                         // cmd_xbar_mux_032:src_valid -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_032_src_startofpacket;                                                                 // cmd_xbar_mux_032:src_startofpacket -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_032_src_data;                                                                          // cmd_xbar_mux_032:src_data -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_032_src_channel;                                                                       // cmd_xbar_mux_032:src_channel -> dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_032_src_ready;                                                                         // dtoe_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_032:src_ready
	wire         id_router_032_src_endofpacket;                                                                      // id_router_032:src_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	wire         id_router_032_src_valid;                                                                            // id_router_032:src_valid -> rsp_xbar_demux_032:sink_valid
	wire         id_router_032_src_startofpacket;                                                                    // id_router_032:src_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	wire  [94:0] id_router_032_src_data;                                                                             // id_router_032:src_data -> rsp_xbar_demux_032:sink_data
	wire  [65:0] id_router_032_src_channel;                                                                          // id_router_032:src_channel -> rsp_xbar_demux_032:sink_channel
	wire         id_router_032_src_ready;                                                                            // rsp_xbar_demux_032:sink_ready -> id_router_032:src_ready
	wire         cmd_xbar_mux_033_src_endofpacket;                                                                   // cmd_xbar_mux_033:src_endofpacket -> dtoe_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_033_src_valid;                                                                         // cmd_xbar_mux_033:src_valid -> dtoe_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_033_src_startofpacket;                                                                 // cmd_xbar_mux_033:src_startofpacket -> dtoe_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_033_src_data;                                                                          // cmd_xbar_mux_033:src_data -> dtoe_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_033_src_channel;                                                                       // cmd_xbar_mux_033:src_channel -> dtoe_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_033_src_ready;                                                                         // dtoe_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_033:src_ready
	wire         id_router_033_src_endofpacket;                                                                      // id_router_033:src_endofpacket -> rsp_xbar_demux_033:sink_endofpacket
	wire         id_router_033_src_valid;                                                                            // id_router_033:src_valid -> rsp_xbar_demux_033:sink_valid
	wire         id_router_033_src_startofpacket;                                                                    // id_router_033:src_startofpacket -> rsp_xbar_demux_033:sink_startofpacket
	wire  [94:0] id_router_033_src_data;                                                                             // id_router_033:src_data -> rsp_xbar_demux_033:sink_data
	wire  [65:0] id_router_033_src_channel;                                                                          // id_router_033:src_channel -> rsp_xbar_demux_033:sink_channel
	wire         id_router_033_src_ready;                                                                            // rsp_xbar_demux_033:sink_ready -> id_router_033:src_ready
	wire         cmd_xbar_demux_004_src10_ready;                                                                     // data_mem_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src10_ready
	wire         id_router_034_src_endofpacket;                                                                      // id_router_034:src_endofpacket -> rsp_xbar_demux_034:sink_endofpacket
	wire         id_router_034_src_valid;                                                                            // id_router_034:src_valid -> rsp_xbar_demux_034:sink_valid
	wire         id_router_034_src_startofpacket;                                                                    // id_router_034:src_startofpacket -> rsp_xbar_demux_034:sink_startofpacket
	wire  [94:0] id_router_034_src_data;                                                                             // id_router_034:src_data -> rsp_xbar_demux_034:sink_data
	wire  [65:0] id_router_034_src_channel;                                                                          // id_router_034:src_channel -> rsp_xbar_demux_034:sink_channel
	wire         id_router_034_src_ready;                                                                            // rsp_xbar_demux_034:sink_ready -> id_router_034:src_ready
	wire         cmd_xbar_demux_004_src11_ready;                                                                     // jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src11_ready
	wire         id_router_035_src_endofpacket;                                                                      // id_router_035:src_endofpacket -> rsp_xbar_demux_035:sink_endofpacket
	wire         id_router_035_src_valid;                                                                            // id_router_035:src_valid -> rsp_xbar_demux_035:sink_valid
	wire         id_router_035_src_startofpacket;                                                                    // id_router_035:src_startofpacket -> rsp_xbar_demux_035:sink_startofpacket
	wire  [94:0] id_router_035_src_data;                                                                             // id_router_035:src_data -> rsp_xbar_demux_035:sink_data
	wire  [65:0] id_router_035_src_channel;                                                                          // id_router_035:src_channel -> rsp_xbar_demux_035:sink_channel
	wire         id_router_035_src_ready;                                                                            // rsp_xbar_demux_035:sink_ready -> id_router_035:src_ready
	wire         cmd_xbar_demux_004_src12_ready;                                                                     // timer_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src12_ready
	wire         id_router_036_src_endofpacket;                                                                      // id_router_036:src_endofpacket -> rsp_xbar_demux_036:sink_endofpacket
	wire         id_router_036_src_valid;                                                                            // id_router_036:src_valid -> rsp_xbar_demux_036:sink_valid
	wire         id_router_036_src_startofpacket;                                                                    // id_router_036:src_startofpacket -> rsp_xbar_demux_036:sink_startofpacket
	wire  [94:0] id_router_036_src_data;                                                                             // id_router_036:src_data -> rsp_xbar_demux_036:sink_data
	wire  [65:0] id_router_036_src_channel;                                                                          // id_router_036:src_channel -> rsp_xbar_demux_036:sink_channel
	wire         id_router_036_src_ready;                                                                            // rsp_xbar_demux_036:sink_ready -> id_router_036:src_ready
	wire         cmd_xbar_demux_004_src13_ready;                                                                     // high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src13_ready
	wire         id_router_037_src_endofpacket;                                                                      // id_router_037:src_endofpacket -> rsp_xbar_demux_037:sink_endofpacket
	wire         id_router_037_src_valid;                                                                            // id_router_037:src_valid -> rsp_xbar_demux_037:sink_valid
	wire         id_router_037_src_startofpacket;                                                                    // id_router_037:src_startofpacket -> rsp_xbar_demux_037:sink_startofpacket
	wire  [94:0] id_router_037_src_data;                                                                             // id_router_037:src_data -> rsp_xbar_demux_037:sink_data
	wire  [65:0] id_router_037_src_channel;                                                                          // id_router_037:src_channel -> rsp_xbar_demux_037:sink_channel
	wire         id_router_037_src_ready;                                                                            // rsp_xbar_demux_037:sink_ready -> id_router_037:src_ready
	wire         cmd_xbar_demux_005_src6_ready;                                                                      // ins_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src6_ready
	wire         id_router_038_src_endofpacket;                                                                      // id_router_038:src_endofpacket -> rsp_xbar_demux_038:sink_endofpacket
	wire         id_router_038_src_valid;                                                                            // id_router_038:src_valid -> rsp_xbar_demux_038:sink_valid
	wire         id_router_038_src_startofpacket;                                                                    // id_router_038:src_startofpacket -> rsp_xbar_demux_038:sink_startofpacket
	wire  [94:0] id_router_038_src_data;                                                                             // id_router_038:src_data -> rsp_xbar_demux_038:sink_data
	wire  [65:0] id_router_038_src_channel;                                                                          // id_router_038:src_channel -> rsp_xbar_demux_038:sink_channel
	wire         id_router_038_src_ready;                                                                            // rsp_xbar_demux_038:sink_ready -> id_router_038:src_ready
	wire         cmd_xbar_mux_039_src_endofpacket;                                                                   // cmd_xbar_mux_039:src_endofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_039_src_valid;                                                                         // cmd_xbar_mux_039:src_valid -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_039_src_startofpacket;                                                                 // cmd_xbar_mux_039:src_startofpacket -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_039_src_data;                                                                          // cmd_xbar_mux_039:src_data -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_039_src_channel;                                                                       // cmd_xbar_mux_039:src_channel -> cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_039_src_ready;                                                                         // cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_039:src_ready
	wire         id_router_039_src_endofpacket;                                                                      // id_router_039:src_endofpacket -> rsp_xbar_demux_039:sink_endofpacket
	wire         id_router_039_src_valid;                                                                            // id_router_039:src_valid -> rsp_xbar_demux_039:sink_valid
	wire         id_router_039_src_startofpacket;                                                                    // id_router_039:src_startofpacket -> rsp_xbar_demux_039:sink_startofpacket
	wire  [94:0] id_router_039_src_data;                                                                             // id_router_039:src_data -> rsp_xbar_demux_039:sink_data
	wire  [65:0] id_router_039_src_channel;                                                                          // id_router_039:src_channel -> rsp_xbar_demux_039:sink_channel
	wire         id_router_039_src_ready;                                                                            // rsp_xbar_demux_039:sink_ready -> id_router_039:src_ready
	wire         cmd_xbar_mux_040_src_endofpacket;                                                                   // cmd_xbar_mux_040:src_endofpacket -> ctod_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_040_src_valid;                                                                         // cmd_xbar_mux_040:src_valid -> ctod_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_040_src_startofpacket;                                                                 // cmd_xbar_mux_040:src_startofpacket -> ctod_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_040_src_data;                                                                          // cmd_xbar_mux_040:src_data -> ctod_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_040_src_channel;                                                                       // cmd_xbar_mux_040:src_channel -> ctod_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_040_src_ready;                                                                         // ctod_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_040:src_ready
	wire         id_router_040_src_endofpacket;                                                                      // id_router_040:src_endofpacket -> rsp_xbar_demux_040:sink_endofpacket
	wire         id_router_040_src_valid;                                                                            // id_router_040:src_valid -> rsp_xbar_demux_040:sink_valid
	wire         id_router_040_src_startofpacket;                                                                    // id_router_040:src_startofpacket -> rsp_xbar_demux_040:sink_startofpacket
	wire  [94:0] id_router_040_src_data;                                                                             // id_router_040:src_data -> rsp_xbar_demux_040:sink_data
	wire  [65:0] id_router_040_src_channel;                                                                          // id_router_040:src_channel -> rsp_xbar_demux_040:sink_channel
	wire         id_router_040_src_ready;                                                                            // rsp_xbar_demux_040:sink_ready -> id_router_040:src_ready
	wire         cmd_xbar_mux_041_src_endofpacket;                                                                   // cmd_xbar_mux_041:src_endofpacket -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_041_src_valid;                                                                         // cmd_xbar_mux_041:src_valid -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_041_src_startofpacket;                                                                 // cmd_xbar_mux_041:src_startofpacket -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_041_src_data;                                                                          // cmd_xbar_mux_041:src_data -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_041_src_channel;                                                                       // cmd_xbar_mux_041:src_channel -> ctod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_041_src_ready;                                                                         // ctod_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_041:src_ready
	wire         id_router_041_src_endofpacket;                                                                      // id_router_041:src_endofpacket -> rsp_xbar_demux_041:sink_endofpacket
	wire         id_router_041_src_valid;                                                                            // id_router_041:src_valid -> rsp_xbar_demux_041:sink_valid
	wire         id_router_041_src_startofpacket;                                                                    // id_router_041:src_startofpacket -> rsp_xbar_demux_041:sink_startofpacket
	wire  [94:0] id_router_041_src_data;                                                                             // id_router_041:src_data -> rsp_xbar_demux_041:sink_data
	wire  [65:0] id_router_041_src_channel;                                                                          // id_router_041:src_channel -> rsp_xbar_demux_041:sink_channel
	wire         id_router_041_src_ready;                                                                            // rsp_xbar_demux_041:sink_ready -> id_router_041:src_ready
	wire         cmd_xbar_mux_042_src_endofpacket;                                                                   // cmd_xbar_mux_042:src_endofpacket -> ctod_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_042_src_valid;                                                                         // cmd_xbar_mux_042:src_valid -> ctod_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_042_src_startofpacket;                                                                 // cmd_xbar_mux_042:src_startofpacket -> ctod_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_042_src_data;                                                                          // cmd_xbar_mux_042:src_data -> ctod_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_042_src_channel;                                                                       // cmd_xbar_mux_042:src_channel -> ctod_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_042_src_ready;                                                                         // ctod_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_042:src_ready
	wire         id_router_042_src_endofpacket;                                                                      // id_router_042:src_endofpacket -> rsp_xbar_demux_042:sink_endofpacket
	wire         id_router_042_src_valid;                                                                            // id_router_042:src_valid -> rsp_xbar_demux_042:sink_valid
	wire         id_router_042_src_startofpacket;                                                                    // id_router_042:src_startofpacket -> rsp_xbar_demux_042:sink_startofpacket
	wire  [94:0] id_router_042_src_data;                                                                             // id_router_042:src_data -> rsp_xbar_demux_042:sink_data
	wire  [65:0] id_router_042_src_channel;                                                                          // id_router_042:src_channel -> rsp_xbar_demux_042:sink_channel
	wire         id_router_042_src_ready;                                                                            // rsp_xbar_demux_042:sink_ready -> id_router_042:src_ready
	wire         cmd_xbar_demux_006_src10_ready;                                                                     // data_mem_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src10_ready
	wire         id_router_043_src_endofpacket;                                                                      // id_router_043:src_endofpacket -> rsp_xbar_demux_043:sink_endofpacket
	wire         id_router_043_src_valid;                                                                            // id_router_043:src_valid -> rsp_xbar_demux_043:sink_valid
	wire         id_router_043_src_startofpacket;                                                                    // id_router_043:src_startofpacket -> rsp_xbar_demux_043:sink_startofpacket
	wire  [94:0] id_router_043_src_data;                                                                             // id_router_043:src_data -> rsp_xbar_demux_043:sink_data
	wire  [65:0] id_router_043_src_channel;                                                                          // id_router_043:src_channel -> rsp_xbar_demux_043:sink_channel
	wire         id_router_043_src_ready;                                                                            // rsp_xbar_demux_043:sink_ready -> id_router_043:src_ready
	wire         cmd_xbar_demux_006_src11_ready;                                                                     // jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src11_ready
	wire         id_router_044_src_endofpacket;                                                                      // id_router_044:src_endofpacket -> rsp_xbar_demux_044:sink_endofpacket
	wire         id_router_044_src_valid;                                                                            // id_router_044:src_valid -> rsp_xbar_demux_044:sink_valid
	wire         id_router_044_src_startofpacket;                                                                    // id_router_044:src_startofpacket -> rsp_xbar_demux_044:sink_startofpacket
	wire  [94:0] id_router_044_src_data;                                                                             // id_router_044:src_data -> rsp_xbar_demux_044:sink_data
	wire  [65:0] id_router_044_src_channel;                                                                          // id_router_044:src_channel -> rsp_xbar_demux_044:sink_channel
	wire         id_router_044_src_ready;                                                                            // rsp_xbar_demux_044:sink_ready -> id_router_044:src_ready
	wire         cmd_xbar_demux_006_src12_ready;                                                                     // timer_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src12_ready
	wire         id_router_045_src_endofpacket;                                                                      // id_router_045:src_endofpacket -> rsp_xbar_demux_045:sink_endofpacket
	wire         id_router_045_src_valid;                                                                            // id_router_045:src_valid -> rsp_xbar_demux_045:sink_valid
	wire         id_router_045_src_startofpacket;                                                                    // id_router_045:src_startofpacket -> rsp_xbar_demux_045:sink_startofpacket
	wire  [94:0] id_router_045_src_data;                                                                             // id_router_045:src_data -> rsp_xbar_demux_045:sink_data
	wire  [65:0] id_router_045_src_channel;                                                                          // id_router_045:src_channel -> rsp_xbar_demux_045:sink_channel
	wire         id_router_045_src_ready;                                                                            // rsp_xbar_demux_045:sink_ready -> id_router_045:src_ready
	wire         cmd_xbar_demux_006_src13_ready;                                                                     // high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_006:src13_ready
	wire         id_router_046_src_endofpacket;                                                                      // id_router_046:src_endofpacket -> rsp_xbar_demux_046:sink_endofpacket
	wire         id_router_046_src_valid;                                                                            // id_router_046:src_valid -> rsp_xbar_demux_046:sink_valid
	wire         id_router_046_src_startofpacket;                                                                    // id_router_046:src_startofpacket -> rsp_xbar_demux_046:sink_startofpacket
	wire  [94:0] id_router_046_src_data;                                                                             // id_router_046:src_data -> rsp_xbar_demux_046:sink_data
	wire  [65:0] id_router_046_src_channel;                                                                          // id_router_046:src_channel -> rsp_xbar_demux_046:sink_channel
	wire         id_router_046_src_ready;                                                                            // rsp_xbar_demux_046:sink_ready -> id_router_046:src_ready
	wire         cmd_xbar_demux_007_src3_ready;                                                                      // data_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src3_ready
	wire         id_router_047_src_endofpacket;                                                                      // id_router_047:src_endofpacket -> rsp_xbar_demux_047:sink_endofpacket
	wire         id_router_047_src_valid;                                                                            // id_router_047:src_valid -> rsp_xbar_demux_047:sink_valid
	wire         id_router_047_src_startofpacket;                                                                    // id_router_047:src_startofpacket -> rsp_xbar_demux_047:sink_startofpacket
	wire  [94:0] id_router_047_src_data;                                                                             // id_router_047:src_data -> rsp_xbar_demux_047:sink_data
	wire  [65:0] id_router_047_src_channel;                                                                          // id_router_047:src_channel -> rsp_xbar_demux_047:sink_channel
	wire         id_router_047_src_ready;                                                                            // rsp_xbar_demux_047:sink_ready -> id_router_047:src_ready
	wire         cmd_xbar_mux_048_src_endofpacket;                                                                   // cmd_xbar_mux_048:src_endofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_048_src_valid;                                                                         // cmd_xbar_mux_048:src_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_048_src_startofpacket;                                                                 // cmd_xbar_mux_048:src_startofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_048_src_data;                                                                          // cmd_xbar_mux_048:src_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_048_src_channel;                                                                       // cmd_xbar_mux_048:src_channel -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_048_src_ready;                                                                         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_048:src_ready
	wire         id_router_048_src_endofpacket;                                                                      // id_router_048:src_endofpacket -> rsp_xbar_demux_048:sink_endofpacket
	wire         id_router_048_src_valid;                                                                            // id_router_048:src_valid -> rsp_xbar_demux_048:sink_valid
	wire         id_router_048_src_startofpacket;                                                                    // id_router_048:src_startofpacket -> rsp_xbar_demux_048:sink_startofpacket
	wire  [94:0] id_router_048_src_data;                                                                             // id_router_048:src_data -> rsp_xbar_demux_048:sink_data
	wire  [65:0] id_router_048_src_channel;                                                                          // id_router_048:src_channel -> rsp_xbar_demux_048:sink_channel
	wire         id_router_048_src_ready;                                                                            // rsp_xbar_demux_048:sink_ready -> id_router_048:src_ready
	wire         cmd_xbar_demux_007_src5_ready;                                                                      // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src5_ready
	wire         id_router_049_src_endofpacket;                                                                      // id_router_049:src_endofpacket -> rsp_xbar_demux_049:sink_endofpacket
	wire         id_router_049_src_valid;                                                                            // id_router_049:src_valid -> rsp_xbar_demux_049:sink_valid
	wire         id_router_049_src_startofpacket;                                                                    // id_router_049:src_startofpacket -> rsp_xbar_demux_049:sink_startofpacket
	wire  [94:0] id_router_049_src_data;                                                                             // id_router_049:src_data -> rsp_xbar_demux_049:sink_data
	wire  [65:0] id_router_049_src_channel;                                                                          // id_router_049:src_channel -> rsp_xbar_demux_049:sink_channel
	wire         id_router_049_src_ready;                                                                            // rsp_xbar_demux_049:sink_ready -> id_router_049:src_ready
	wire         cmd_xbar_demux_007_src6_ready;                                                                      // timer_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src6_ready
	wire         id_router_050_src_endofpacket;                                                                      // id_router_050:src_endofpacket -> rsp_xbar_demux_050:sink_endofpacket
	wire         id_router_050_src_valid;                                                                            // id_router_050:src_valid -> rsp_xbar_demux_050:sink_valid
	wire         id_router_050_src_startofpacket;                                                                    // id_router_050:src_startofpacket -> rsp_xbar_demux_050:sink_startofpacket
	wire  [94:0] id_router_050_src_data;                                                                             // id_router_050:src_data -> rsp_xbar_demux_050:sink_data
	wire  [65:0] id_router_050_src_channel;                                                                          // id_router_050:src_channel -> rsp_xbar_demux_050:sink_channel
	wire         id_router_050_src_ready;                                                                            // rsp_xbar_demux_050:sink_ready -> id_router_050:src_ready
	wire         cmd_xbar_demux_007_src7_ready;                                                                      // high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src7_ready
	wire         id_router_051_src_endofpacket;                                                                      // id_router_051:src_endofpacket -> rsp_xbar_demux_051:sink_endofpacket
	wire         id_router_051_src_valid;                                                                            // id_router_051:src_valid -> rsp_xbar_demux_051:sink_valid
	wire         id_router_051_src_startofpacket;                                                                    // id_router_051:src_startofpacket -> rsp_xbar_demux_051:sink_startofpacket
	wire  [94:0] id_router_051_src_data;                                                                             // id_router_051:src_data -> rsp_xbar_demux_051:sink_data
	wire  [65:0] id_router_051_src_channel;                                                                          // id_router_051:src_channel -> rsp_xbar_demux_051:sink_channel
	wire         id_router_051_src_ready;                                                                            // rsp_xbar_demux_051:sink_ready -> id_router_051:src_ready
	wire         cmd_xbar_mux_052_src_endofpacket;                                                                   // cmd_xbar_mux_052:src_endofpacket -> btoc_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_052_src_valid;                                                                         // cmd_xbar_mux_052:src_valid -> btoc_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_052_src_startofpacket;                                                                 // cmd_xbar_mux_052:src_startofpacket -> btoc_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_052_src_data;                                                                          // cmd_xbar_mux_052:src_data -> btoc_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_052_src_channel;                                                                       // cmd_xbar_mux_052:src_channel -> btoc_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_052_src_ready;                                                                         // btoc_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_052:src_ready
	wire         id_router_052_src_endofpacket;                                                                      // id_router_052:src_endofpacket -> rsp_xbar_demux_052:sink_endofpacket
	wire         id_router_052_src_valid;                                                                            // id_router_052:src_valid -> rsp_xbar_demux_052:sink_valid
	wire         id_router_052_src_startofpacket;                                                                    // id_router_052:src_startofpacket -> rsp_xbar_demux_052:sink_startofpacket
	wire  [94:0] id_router_052_src_data;                                                                             // id_router_052:src_data -> rsp_xbar_demux_052:sink_data
	wire  [65:0] id_router_052_src_channel;                                                                          // id_router_052:src_channel -> rsp_xbar_demux_052:sink_channel
	wire         id_router_052_src_ready;                                                                            // rsp_xbar_demux_052:sink_ready -> id_router_052:src_ready
	wire         cmd_xbar_mux_053_src_endofpacket;                                                                   // cmd_xbar_mux_053:src_endofpacket -> btoc_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_053_src_valid;                                                                         // cmd_xbar_mux_053:src_valid -> btoc_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_053_src_startofpacket;                                                                 // cmd_xbar_mux_053:src_startofpacket -> btoc_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_053_src_data;                                                                          // cmd_xbar_mux_053:src_data -> btoc_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_053_src_channel;                                                                       // cmd_xbar_mux_053:src_channel -> btoc_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_053_src_ready;                                                                         // btoc_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_053:src_ready
	wire         id_router_053_src_endofpacket;                                                                      // id_router_053:src_endofpacket -> rsp_xbar_demux_053:sink_endofpacket
	wire         id_router_053_src_valid;                                                                            // id_router_053:src_valid -> rsp_xbar_demux_053:sink_valid
	wire         id_router_053_src_startofpacket;                                                                    // id_router_053:src_startofpacket -> rsp_xbar_demux_053:sink_startofpacket
	wire  [94:0] id_router_053_src_data;                                                                             // id_router_053:src_data -> rsp_xbar_demux_053:sink_data
	wire  [65:0] id_router_053_src_channel;                                                                          // id_router_053:src_channel -> rsp_xbar_demux_053:sink_channel
	wire         id_router_053_src_ready;                                                                            // rsp_xbar_demux_053:sink_ready -> id_router_053:src_ready
	wire         cmd_xbar_mux_054_src_endofpacket;                                                                   // cmd_xbar_mux_054:src_endofpacket -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_054_src_valid;                                                                         // cmd_xbar_mux_054:src_valid -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_054_src_startofpacket;                                                                 // cmd_xbar_mux_054:src_startofpacket -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_054_src_data;                                                                          // cmd_xbar_mux_054:src_data -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_054_src_channel;                                                                       // cmd_xbar_mux_054:src_channel -> btoc_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_054_src_ready;                                                                         // btoc_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_054:src_ready
	wire         id_router_054_src_endofpacket;                                                                      // id_router_054:src_endofpacket -> rsp_xbar_demux_054:sink_endofpacket
	wire         id_router_054_src_valid;                                                                            // id_router_054:src_valid -> rsp_xbar_demux_054:sink_valid
	wire         id_router_054_src_startofpacket;                                                                    // id_router_054:src_startofpacket -> rsp_xbar_demux_054:sink_startofpacket
	wire  [94:0] id_router_054_src_data;                                                                             // id_router_054:src_data -> rsp_xbar_demux_054:sink_data
	wire  [65:0] id_router_054_src_channel;                                                                          // id_router_054:src_channel -> rsp_xbar_demux_054:sink_channel
	wire         id_router_054_src_ready;                                                                            // rsp_xbar_demux_054:sink_ready -> id_router_054:src_ready
	wire         cmd_xbar_demux_008_src7_ready;                                                                      // ins_mem_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src7_ready
	wire         id_router_055_src_endofpacket;                                                                      // id_router_055:src_endofpacket -> rsp_xbar_demux_055:sink_endofpacket
	wire         id_router_055_src_valid;                                                                            // id_router_055:src_valid -> rsp_xbar_demux_055:sink_valid
	wire         id_router_055_src_startofpacket;                                                                    // id_router_055:src_startofpacket -> rsp_xbar_demux_055:sink_startofpacket
	wire  [94:0] id_router_055_src_data;                                                                             // id_router_055:src_data -> rsp_xbar_demux_055:sink_data
	wire  [65:0] id_router_055_src_channel;                                                                          // id_router_055:src_channel -> rsp_xbar_demux_055:sink_channel
	wire         id_router_055_src_ready;                                                                            // rsp_xbar_demux_055:sink_ready -> id_router_055:src_ready
	wire         cmd_xbar_demux_009_src12_ready;                                                                     // ins_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_009:src12_ready
	wire         id_router_056_src_endofpacket;                                                                      // id_router_056:src_endofpacket -> rsp_xbar_demux_056:sink_endofpacket
	wire         id_router_056_src_valid;                                                                            // id_router_056:src_valid -> rsp_xbar_demux_056:sink_valid
	wire         id_router_056_src_startofpacket;                                                                    // id_router_056:src_startofpacket -> rsp_xbar_demux_056:sink_startofpacket
	wire  [94:0] id_router_056_src_data;                                                                             // id_router_056:src_data -> rsp_xbar_demux_056:sink_data
	wire  [65:0] id_router_056_src_channel;                                                                          // id_router_056:src_channel -> rsp_xbar_demux_056:sink_channel
	wire         id_router_056_src_ready;                                                                            // rsp_xbar_demux_056:sink_ready -> id_router_056:src_ready
	wire         cmd_xbar_mux_057_src_endofpacket;                                                                   // cmd_xbar_mux_057:src_endofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_057_src_valid;                                                                         // cmd_xbar_mux_057:src_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_057_src_startofpacket;                                                                 // cmd_xbar_mux_057:src_startofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_057_src_data;                                                                          // cmd_xbar_mux_057:src_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [65:0] cmd_xbar_mux_057_src_channel;                                                                       // cmd_xbar_mux_057:src_channel -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_057_src_ready;                                                                         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_057:src_ready
	wire         id_router_057_src_endofpacket;                                                                      // id_router_057:src_endofpacket -> rsp_xbar_demux_057:sink_endofpacket
	wire         id_router_057_src_valid;                                                                            // id_router_057:src_valid -> rsp_xbar_demux_057:sink_valid
	wire         id_router_057_src_startofpacket;                                                                    // id_router_057:src_startofpacket -> rsp_xbar_demux_057:sink_startofpacket
	wire  [94:0] id_router_057_src_data;                                                                             // id_router_057:src_data -> rsp_xbar_demux_057:sink_data
	wire  [65:0] id_router_057_src_channel;                                                                          // id_router_057:src_channel -> rsp_xbar_demux_057:sink_channel
	wire         id_router_057_src_ready;                                                                            // rsp_xbar_demux_057:sink_ready -> id_router_057:src_ready
	wire         cmd_xbar_demux_010_src13_ready;                                                                     // data_mem_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_010:src13_ready
	wire         id_router_058_src_endofpacket;                                                                      // id_router_058:src_endofpacket -> rsp_xbar_demux_058:sink_endofpacket
	wire         id_router_058_src_valid;                                                                            // id_router_058:src_valid -> rsp_xbar_demux_058:sink_valid
	wire         id_router_058_src_startofpacket;                                                                    // id_router_058:src_startofpacket -> rsp_xbar_demux_058:sink_startofpacket
	wire  [94:0] id_router_058_src_data;                                                                             // id_router_058:src_data -> rsp_xbar_demux_058:sink_data
	wire  [65:0] id_router_058_src_channel;                                                                          // id_router_058:src_channel -> rsp_xbar_demux_058:sink_channel
	wire         id_router_058_src_ready;                                                                            // rsp_xbar_demux_058:sink_ready -> id_router_058:src_ready
	wire         cmd_xbar_demux_010_src14_ready;                                                                     // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_010:src14_ready
	wire         id_router_059_src_endofpacket;                                                                      // id_router_059:src_endofpacket -> rsp_xbar_demux_059:sink_endofpacket
	wire         id_router_059_src_valid;                                                                            // id_router_059:src_valid -> rsp_xbar_demux_059:sink_valid
	wire         id_router_059_src_startofpacket;                                                                    // id_router_059:src_startofpacket -> rsp_xbar_demux_059:sink_startofpacket
	wire  [94:0] id_router_059_src_data;                                                                             // id_router_059:src_data -> rsp_xbar_demux_059:sink_data
	wire  [65:0] id_router_059_src_channel;                                                                          // id_router_059:src_channel -> rsp_xbar_demux_059:sink_channel
	wire         id_router_059_src_ready;                                                                            // rsp_xbar_demux_059:sink_ready -> id_router_059:src_ready
	wire         cmd_xbar_demux_010_src15_ready;                                                                     // timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_010:src15_ready
	wire         id_router_060_src_endofpacket;                                                                      // id_router_060:src_endofpacket -> rsp_xbar_demux_060:sink_endofpacket
	wire         id_router_060_src_valid;                                                                            // id_router_060:src_valid -> rsp_xbar_demux_060:sink_valid
	wire         id_router_060_src_startofpacket;                                                                    // id_router_060:src_startofpacket -> rsp_xbar_demux_060:sink_startofpacket
	wire  [94:0] id_router_060_src_data;                                                                             // id_router_060:src_data -> rsp_xbar_demux_060:sink_data
	wire  [65:0] id_router_060_src_channel;                                                                          // id_router_060:src_channel -> rsp_xbar_demux_060:sink_channel
	wire         id_router_060_src_ready;                                                                            // rsp_xbar_demux_060:sink_ready -> id_router_060:src_ready
	wire         cmd_xbar_demux_010_src16_ready;                                                                     // high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_010:src16_ready
	wire         id_router_061_src_endofpacket;                                                                      // id_router_061:src_endofpacket -> rsp_xbar_demux_061:sink_endofpacket
	wire         id_router_061_src_valid;                                                                            // id_router_061:src_valid -> rsp_xbar_demux_061:sink_valid
	wire         id_router_061_src_startofpacket;                                                                    // id_router_061:src_startofpacket -> rsp_xbar_demux_061:sink_startofpacket
	wire  [94:0] id_router_061_src_data;                                                                             // id_router_061:src_data -> rsp_xbar_demux_061:sink_data
	wire  [65:0] id_router_061_src_channel;                                                                          // id_router_061:src_channel -> rsp_xbar_demux_061:sink_channel
	wire         id_router_061_src_ready;                                                                            // rsp_xbar_demux_061:sink_ready -> id_router_061:src_ready
	wire         cmd_xbar_demux_011_src19_ready;                                                                     // data_mem_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_011:src19_ready
	wire         id_router_062_src_endofpacket;                                                                      // id_router_062:src_endofpacket -> rsp_xbar_demux_062:sink_endofpacket
	wire         id_router_062_src_valid;                                                                            // id_router_062:src_valid -> rsp_xbar_demux_062:sink_valid
	wire         id_router_062_src_startofpacket;                                                                    // id_router_062:src_startofpacket -> rsp_xbar_demux_062:sink_startofpacket
	wire  [94:0] id_router_062_src_data;                                                                             // id_router_062:src_data -> rsp_xbar_demux_062:sink_data
	wire  [65:0] id_router_062_src_channel;                                                                          // id_router_062:src_channel -> rsp_xbar_demux_062:sink_channel
	wire         id_router_062_src_ready;                                                                            // rsp_xbar_demux_062:sink_ready -> id_router_062:src_ready
	wire         cmd_xbar_demux_011_src20_ready;                                                                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_011:src20_ready
	wire         id_router_063_src_endofpacket;                                                                      // id_router_063:src_endofpacket -> rsp_xbar_demux_063:sink_endofpacket
	wire         id_router_063_src_valid;                                                                            // id_router_063:src_valid -> rsp_xbar_demux_063:sink_valid
	wire         id_router_063_src_startofpacket;                                                                    // id_router_063:src_startofpacket -> rsp_xbar_demux_063:sink_startofpacket
	wire  [94:0] id_router_063_src_data;                                                                             // id_router_063:src_data -> rsp_xbar_demux_063:sink_data
	wire  [65:0] id_router_063_src_channel;                                                                          // id_router_063:src_channel -> rsp_xbar_demux_063:sink_channel
	wire         id_router_063_src_ready;                                                                            // rsp_xbar_demux_063:sink_ready -> id_router_063:src_ready
	wire         cmd_xbar_demux_011_src21_ready;                                                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_011:src21_ready
	wire         id_router_064_src_endofpacket;                                                                      // id_router_064:src_endofpacket -> rsp_xbar_demux_064:sink_endofpacket
	wire         id_router_064_src_valid;                                                                            // id_router_064:src_valid -> rsp_xbar_demux_064:sink_valid
	wire         id_router_064_src_startofpacket;                                                                    // id_router_064:src_startofpacket -> rsp_xbar_demux_064:sink_startofpacket
	wire  [94:0] id_router_064_src_data;                                                                             // id_router_064:src_data -> rsp_xbar_demux_064:sink_data
	wire  [65:0] id_router_064_src_channel;                                                                          // id_router_064:src_channel -> rsp_xbar_demux_064:sink_channel
	wire         id_router_064_src_ready;                                                                            // rsp_xbar_demux_064:sink_ready -> id_router_064:src_ready
	wire         cmd_xbar_demux_011_src22_ready;                                                                     // high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_011:src22_ready
	wire         id_router_065_src_endofpacket;                                                                      // id_router_065:src_endofpacket -> rsp_xbar_demux_065:sink_endofpacket
	wire         id_router_065_src_valid;                                                                            // id_router_065:src_valid -> rsp_xbar_demux_065:sink_valid
	wire         id_router_065_src_startofpacket;                                                                    // id_router_065:src_startofpacket -> rsp_xbar_demux_065:sink_startofpacket
	wire  [94:0] id_router_065_src_data;                                                                             // id_router_065:src_data -> rsp_xbar_demux_065:sink_data
	wire  [65:0] id_router_065_src_channel;                                                                          // id_router_065:src_channel -> rsp_xbar_demux_065:sink_channel
	wire         id_router_065_src_ready;                                                                            // rsp_xbar_demux_065:sink_ready -> id_router_065:src_ready
	wire  [65:0] limiter_cmd_valid_data;                                                                             // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire  [65:0] limiter_001_cmd_valid_data;                                                                         // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire  [65:0] limiter_002_cmd_valid_data;                                                                         // limiter_002:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire  [65:0] limiter_003_cmd_valid_data;                                                                         // limiter_003:cmd_src_valid -> cmd_xbar_demux_005:sink_valid
	wire  [65:0] limiter_004_cmd_valid_data;                                                                         // limiter_004:cmd_src_valid -> cmd_xbar_demux_008:sink_valid
	wire  [65:0] limiter_005_cmd_valid_data;                                                                         // limiter_005:cmd_src_valid -> cmd_xbar_demux_009:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                           // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                           // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                           // high_scale_timer_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_0_d_irq_irq;                                                                                    // irq_mapper:sender_irq -> cpu_0:d_irq
	wire         irq_mapper_001_receiver0_irq;                                                                       // jtag_uart_1:av_irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                                                       // timer_1:irq -> irq_mapper_001:receiver1_irq
	wire         irq_mapper_001_receiver2_irq;                                                                       // high_scale_timer_1:irq -> irq_mapper_001:receiver2_irq
	wire  [31:0] cpu_1_d_irq_irq;                                                                                    // irq_mapper_001:sender_irq -> cpu_1:d_irq
	wire         irq_mapper_002_receiver0_irq;                                                                       // jtag_uart_2:av_irq -> irq_mapper_002:receiver0_irq
	wire         irq_mapper_002_receiver1_irq;                                                                       // timer_2:irq -> irq_mapper_002:receiver1_irq
	wire         irq_mapper_002_receiver2_irq;                                                                       // high_scale_timer_2:irq -> irq_mapper_002:receiver2_irq
	wire  [31:0] cpu_2_d_irq_irq;                                                                                    // irq_mapper_002:sender_irq -> cpu_2:d_irq
	wire         irq_mapper_003_receiver0_irq;                                                                       // jtag_uart_3:av_irq -> irq_mapper_003:receiver0_irq
	wire         irq_mapper_003_receiver1_irq;                                                                       // timer_3:irq -> irq_mapper_003:receiver1_irq
	wire         irq_mapper_003_receiver2_irq;                                                                       // high_scale_timer_3:irq -> irq_mapper_003:receiver2_irq
	wire  [31:0] cpu_3_d_irq_irq;                                                                                    // irq_mapper_003:sender_irq -> cpu_3:d_irq
	wire         irq_mapper_004_receiver0_irq;                                                                       // jtag_uart_4:av_irq -> irq_mapper_004:receiver0_irq
	wire         irq_mapper_004_receiver1_irq;                                                                       // timer_4:irq -> irq_mapper_004:receiver1_irq
	wire         irq_mapper_004_receiver2_irq;                                                                       // high_scale_timer_4:irq -> irq_mapper_004:receiver2_irq
	wire  [31:0] cpu_4_d_irq_irq;                                                                                    // irq_mapper_004:sender_irq -> cpu_4:d_irq
	wire         irq_mapper_005_receiver0_irq;                                                                       // jtag_uart_5:av_irq -> irq_mapper_005:receiver0_irq
	wire         irq_mapper_005_receiver1_irq;                                                                       // timer_5:irq -> irq_mapper_005:receiver1_irq
	wire         irq_mapper_005_receiver2_irq;                                                                       // high_scale_timer_5:irq -> irq_mapper_005:receiver2_irq
	wire  [31:0] cpu_5_d_irq_irq;                                                                                    // irq_mapper_005:sender_irq -> cpu_5:d_irq
	wire         irq_mapper_receiver3_irq;                                                                           // atob_0:wrclk_control_slave_irq -> [irq_mapper:receiver3_irq, irq_mapper_001:receiver3_irq]
	wire         irq_mapper_receiver4_irq;                                                                           // atob_1:wrclk_control_slave_irq -> [irq_mapper:receiver4_irq, irq_mapper_001:receiver4_irq]
	wire         irq_mapper_receiver5_irq;                                                                           // atob_2:wrclk_control_slave_irq -> [irq_mapper:receiver5_irq, irq_mapper_001:receiver5_irq]
	wire         irq_mapper_001_receiver6_irq;                                                                       // btoc_0:wrclk_control_slave_irq -> [irq_mapper_001:receiver6_irq, irq_mapper_002:receiver3_irq]
	wire         irq_mapper_002_receiver4_irq;                                                                       // ctod_0:wrclk_control_slave_irq -> [irq_mapper_002:receiver4_irq, irq_mapper_003:receiver3_irq]
	wire         irq_mapper_003_receiver4_irq;                                                                       // dtoe_0:wrclk_control_slave_irq -> [irq_mapper_003:receiver4_irq, irq_mapper_004:receiver3_irq]
	wire         irq_mapper_004_receiver4_irq;                                                                       // etof_0:wrclk_control_slave_irq -> [irq_mapper_004:receiver4_irq, irq_mapper_005:receiver3_irq]
	wire         irq_mapper_receiver8_irq;                                                                           // atof_0:wrclk_control_slave_irq -> [irq_mapper:receiver8_irq, irq_mapper_005:receiver4_irq]
	wire         irq_mapper_receiver6_irq;                                                                           // atod_0:wrclk_control_slave_irq -> [irq_mapper:receiver6_irq, irq_mapper_003:receiver5_irq]
	wire         irq_mapper_receiver7_irq;                                                                           // atoe_0:wrclk_control_slave_irq -> [irq_mapper:receiver7_irq, irq_mapper_004:receiver5_irq]

	SoC_ins_mem_0 ins_mem_0 (
		.clk        (clk_clk),                                                //   clk1.clk
		.address    (ins_mem_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ins_mem_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ins_mem_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ins_mem_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ins_mem_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ins_mem_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ins_mem_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                          // reset1.reset
	);

	SoC_data_mem_0 data_mem_0 (
		.clk        (clk_clk),                                                 //   clk1.clk
		.address    (data_mem_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (data_mem_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (data_mem_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (data_mem_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (data_mem_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (data_mem_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (data_mem_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                           // reset1.reset
	);

	SoC_cpu_0 cpu_0 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (cpu_0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_0_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_0_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_0_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_0_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                  //               irq.irq
	);

	SoC_timer_0 timer_0 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                              //   irq.irq
	);

	SoC_high_scale_timer_0 high_scale_timer_0 (
		.clk        (clk_clk),                                                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                 // reset.reset_n
		.address    (high_scale_timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_scale_timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_scale_timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_scale_timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_scale_timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                                         //   irq.irq
	);

	SoC_ins_mem_1 ins_mem_1 (
		.clk        (clk_clk),                                                //   clk1.clk
		.address    (ins_mem_1_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ins_mem_1_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ins_mem_1_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ins_mem_1_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ins_mem_1_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ins_mem_1_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ins_mem_1_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset)                      // reset1.reset
	);

	SoC_data_mem_1 data_mem_1 (
		.clk        (clk_clk),                                                 //   clk1.clk
		.address    (data_mem_1_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (data_mem_1_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (data_mem_1_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (data_mem_1_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (data_mem_1_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (data_mem_1_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (data_mem_1_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset)                       // reset1.reset
	);

	SoC_cpu_1 cpu_1 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                                  //                   reset_n.reset_n
		.d_address                             (cpu_1_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_1_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_1_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_1_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_1_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_1_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_1_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_1_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_1_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_1_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_1_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_1_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_1_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_1 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver0_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_1 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  // reset.reset_n
		.address    (timer_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_001_receiver1_irq)                          //   irq.irq
	);

	SoC_high_scale_timer_0 high_scale_timer_1 (
		.clk        (clk_clk),                                                         //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                             // reset.reset_n
		.address    (high_scale_timer_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_scale_timer_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_scale_timer_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_scale_timer_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_scale_timer_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_001_receiver2_irq)                                     //   irq.irq
	);

	SoC_ins_mem_2 ins_mem_2 (
		.clk        (clk_clk),                                                //   clk1.clk
		.address    (ins_mem_2_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ins_mem_2_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ins_mem_2_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ins_mem_2_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ins_mem_2_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ins_mem_2_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ins_mem_2_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset)                      // reset1.reset
	);

	SoC_data_mem_2 data_mem_2 (
		.clk        (clk_clk),                                                 //   clk1.clk
		.address    (data_mem_2_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (data_mem_2_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (data_mem_2_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (data_mem_2_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (data_mem_2_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (data_mem_2_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (data_mem_2_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset)                       // reset1.reset
	);

	SoC_cpu_2 cpu_2 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_003_reset_out_reset),                                  //                   reset_n.reset_n
		.d_address                             (cpu_2_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_2_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_2_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_2_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_2_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_2_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_2_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_2_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_2_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_2_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_2_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_2_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_2_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_2_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_2_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_2 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver0_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_2 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                  // reset.reset_n
		.address    (timer_2_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_2_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_2_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_2_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_2_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_002_receiver1_irq)                          //   irq.irq
	);

	SoC_high_scale_timer_0 high_scale_timer_2 (
		.clk        (clk_clk),                                                         //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                             // reset.reset_n
		.address    (high_scale_timer_2_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_scale_timer_2_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_scale_timer_2_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_scale_timer_2_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_scale_timer_2_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_002_receiver2_irq)                                     //   irq.irq
	);

	SoC_ins_mem_3 ins_mem_3 (
		.clk        (clk_clk),                                                //   clk1.clk
		.address    (ins_mem_3_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ins_mem_3_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ins_mem_3_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ins_mem_3_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ins_mem_3_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ins_mem_3_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ins_mem_3_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_004_reset_out_reset)                      // reset1.reset
	);

	SoC_data_mem_3 data_mem_3 (
		.clk        (clk_clk),                                                 //   clk1.clk
		.address    (data_mem_3_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (data_mem_3_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (data_mem_3_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (data_mem_3_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (data_mem_3_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (data_mem_3_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (data_mem_3_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_004_reset_out_reset)                       // reset1.reset
	);

	SoC_cpu_3 cpu_3 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_004_reset_out_reset),                                  //                   reset_n.reset_n
		.d_address                             (cpu_3_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_3_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_3_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_3_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_3_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_3_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_3_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_3_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_3_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_3_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_3_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_3_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_3_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_3_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_3_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_3 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_004_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_003_receiver0_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_3 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                  // reset.reset_n
		.address    (timer_3_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_3_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_3_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_3_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_3_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_003_receiver1_irq)                          //   irq.irq
	);

	SoC_high_scale_timer_0 high_scale_timer_3 (
		.clk        (clk_clk),                                                         //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                             // reset.reset_n
		.address    (high_scale_timer_3_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_scale_timer_3_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_scale_timer_3_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_scale_timer_3_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_scale_timer_3_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_003_receiver2_irq)                                     //   irq.irq
	);

	SoC_ins_mem_4 ins_mem_4 (
		.clk        (clk_clk),                                                //   clk1.clk
		.address    (ins_mem_4_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ins_mem_4_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ins_mem_4_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ins_mem_4_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ins_mem_4_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ins_mem_4_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ins_mem_4_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_005_reset_out_reset)                      // reset1.reset
	);

	SoC_data_mem_4 data_mem_4 (
		.clk        (clk_clk),                                                 //   clk1.clk
		.address    (data_mem_4_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (data_mem_4_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (data_mem_4_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (data_mem_4_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (data_mem_4_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (data_mem_4_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (data_mem_4_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_005_reset_out_reset)                       // reset1.reset
	);

	SoC_cpu_4 cpu_4 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_005_reset_out_reset),                                  //                   reset_n.reset_n
		.d_address                             (cpu_4_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_4_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_4_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_4_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_4_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_4_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_4_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_4_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_4_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_4_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_4_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_4_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_4_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_4_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_4_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_4 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_005_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_004_receiver0_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_4 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_005_reset_out_reset),                  // reset.reset_n
		.address    (timer_4_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_4_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_4_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_4_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_4_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_004_receiver1_irq)                          //   irq.irq
	);

	SoC_high_scale_timer_0 high_scale_timer_4 (
		.clk        (clk_clk),                                                         //   clk.clk
		.reset_n    (~rst_controller_005_reset_out_reset),                             // reset.reset_n
		.address    (high_scale_timer_4_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_scale_timer_4_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_scale_timer_4_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_scale_timer_4_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_scale_timer_4_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_004_receiver2_irq)                                     //   irq.irq
	);

	SoC_ins_mem_5 ins_mem_5 (
		.clk        (clk_clk),                                                //   clk1.clk
		.address    (ins_mem_5_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ins_mem_5_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ins_mem_5_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ins_mem_5_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ins_mem_5_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ins_mem_5_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ins_mem_5_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_006_reset_out_reset)                      // reset1.reset
	);

	SoC_data_mem_5 data_mem_5 (
		.clk        (clk_clk),                                                 //   clk1.clk
		.address    (data_mem_5_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (data_mem_5_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (data_mem_5_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (data_mem_5_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (data_mem_5_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (data_mem_5_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (data_mem_5_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_006_reset_out_reset)                       // reset1.reset
	);

	SoC_cpu_5 cpu_5 (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_006_reset_out_reset),                                  //                   reset_n.reset_n
		.d_address                             (cpu_5_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_5_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_5_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_5_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_5_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_5_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_5_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_5_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_5_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_5_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_5_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_5_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_5_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_5_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_5_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SoC_jtag_uart_0 jtag_uart_5 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_006_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_005_receiver0_irq)                                              //               irq.irq
	);

	SoC_timer_0 timer_5 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),                  // reset.reset_n
		.address    (timer_5_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_5_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_5_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_5_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_5_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_005_receiver1_irq)                          //   irq.irq
	);

	SoC_high_scale_timer_0 high_scale_timer_5 (
		.clk        (clk_clk),                                                         //   clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),                             // reset.reset_n
		.address    (high_scale_timer_5_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_scale_timer_5_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_scale_timer_5_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_scale_timer_5_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_scale_timer_5_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_005_receiver2_irq)                                     //   irq.irq
	);

	SoC_atob_0 atob_0 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_007_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (atob_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (atob_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (atob_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (atob_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (atob_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (atob_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (atob_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (atob_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver3_irq),                               //   in_irq.irq
		.avalonmm_read_slave_readdata     (atob_0_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (atob_0_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (atob_0_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_atob_0 atob_1 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_007_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (atob_1_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (atob_1_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (atob_1_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (atob_1_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (atob_1_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (atob_1_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (atob_1_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (atob_1_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver4_irq),                               //   in_irq.irq
		.avalonmm_read_slave_readdata     (atob_1_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (atob_1_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (atob_1_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_atob_0 atob_2 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_007_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (atob_2_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (atob_2_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (atob_2_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (atob_2_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (atob_2_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (atob_2_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (atob_2_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (atob_2_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver5_irq),                               //   in_irq.irq
		.avalonmm_read_slave_readdata     (atob_2_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (atob_2_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (atob_2_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_atob_0 btoc_0 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_008_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (btoc_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (btoc_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (btoc_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (btoc_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (btoc_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (btoc_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (btoc_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (btoc_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_001_receiver6_irq),                           //   in_irq.irq
		.avalonmm_read_slave_readdata     (btoc_0_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (btoc_0_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (btoc_0_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_atob_0 ctod_0 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_009_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (ctod_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (ctod_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (ctod_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (ctod_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (ctod_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (ctod_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (ctod_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (ctod_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_002_receiver4_irq),                           //   in_irq.irq
		.avalonmm_read_slave_readdata     (ctod_0_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (ctod_0_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (ctod_0_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_atob_0 dtoe_0 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_010_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (dtoe_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (dtoe_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (dtoe_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (dtoe_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (dtoe_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (dtoe_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (dtoe_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (dtoe_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_003_receiver4_irq),                           //   in_irq.irq
		.avalonmm_read_slave_readdata     (dtoe_0_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (dtoe_0_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (dtoe_0_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_atob_0 etof_0 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_011_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (etof_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (etof_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (etof_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (etof_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (etof_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (etof_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (etof_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (etof_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_004_receiver4_irq),                           //   in_irq.irq
		.avalonmm_read_slave_readdata     (etof_0_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (etof_0_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (etof_0_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_atob_0 atof_0 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_012_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (atof_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (atof_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (atof_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (atof_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (atof_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (atof_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (atof_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (atof_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver8_irq),                               //   in_irq.irq
		.avalonmm_read_slave_readdata     (atof_0_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (atof_0_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (atof_0_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_atob_0 atod_0 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_013_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (atod_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (atod_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (atod_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (atod_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (atod_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (atod_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (atod_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (atod_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver6_irq),                               //   in_irq.irq
		.avalonmm_read_slave_readdata     (atod_0_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (atod_0_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (atod_0_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	SoC_atob_0 atoe_0 (
		.wrclock                          (clk_clk),                                                //   clk_in.clk
		.reset_n                          (~rst_controller_014_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (atoe_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (atoe_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_waitrequest (atoe_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (atoe_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (atoe_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (atoe_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (atoe_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (atoe_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver7_irq),                               //   in_irq.irq
		.avalonmm_read_slave_readdata     (atoe_0_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (atoe_0_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_waitrequest  (atoe_0_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_0_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_0_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_0_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_0_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_5_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                          //                     reset.reset
		.uav_address           (cpu_5_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_5_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_5_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_5_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_5_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_5_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_5_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_5_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_5_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_5_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_5_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_5_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_5_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_5_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_5_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_5_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_5_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                   //                     reset.reset
		.uav_address           (cpu_5_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_5_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_5_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_5_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_5_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_5_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_5_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_5_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_5_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_5_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_5_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_5_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_5_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_5_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_5_data_master_read),                                               //                          .read
		.av_readdata           (cpu_5_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_5_data_master_write),                                              //                          .write
		.av_writedata          (cpu_5_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_5_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_0_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_0_data_master_read),                                               //                          .read
		.av_readdata           (cpu_0_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_0_data_master_write),                                              //                          .write
		.av_writedata          (cpu_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_4_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                          //                     reset.reset
		.uav_address           (cpu_4_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_4_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_4_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_4_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_4_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_4_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_4_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_4_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_4_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_4_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_4_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_4_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_4_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_4_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_4_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_4_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_4_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                   //                     reset.reset
		.uav_address           (cpu_4_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_4_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_4_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_4_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_4_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_4_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_4_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_4_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_4_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_4_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_4_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_4_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_4_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_4_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_4_data_master_read),                                               //                          .read
		.av_readdata           (cpu_4_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_4_data_master_write),                                              //                          .write
		.av_writedata          (cpu_4_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_4_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_3_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                          //                     reset.reset
		.uav_address           (cpu_3_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_3_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_3_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_3_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_3_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_3_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_3_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_3_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_3_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_3_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_3_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_3_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_3_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_3_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_3_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_3_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_3_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                   //                     reset.reset
		.uav_address           (cpu_3_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_3_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_3_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_3_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_3_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_3_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_3_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_3_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_3_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_3_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_3_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_3_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_3_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_3_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_3_data_master_read),                                               //                          .read
		.av_readdata           (cpu_3_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_3_data_master_write),                                              //                          .write
		.av_writedata          (cpu_3_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_3_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_2_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                   //                     reset.reset
		.uav_address           (cpu_2_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_2_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_2_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_2_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_2_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_2_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_2_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_2_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_2_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_2_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_2_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_2_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_2_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_2_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_2_data_master_read),                                               //                          .read
		.av_readdata           (cpu_2_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_2_data_master_write),                                              //                          .write
		.av_writedata          (cpu_2_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_2_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_2_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                          //                     reset.reset
		.uav_address           (cpu_2_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_2_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_2_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_2_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_2_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_2_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_2_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_2_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_2_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_2_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_2_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_2_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_2_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_2_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_2_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_2_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_1_instruction_master_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                          //                     reset.reset
		.uav_address           (cpu_1_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_1_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_1_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_1_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_1_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_1_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_1_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_1_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_1_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_1_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_1_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_1_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_1_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_1_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_1_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_1_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (14),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (14),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_1_data_master_translator (
		.clk                   (clk_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                   //                     reset.reset
		.uav_address           (cpu_1_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_1_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_1_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_1_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_1_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_1_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_1_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_1_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_1_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_1_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_1_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_1_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_1_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_1_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_1_data_master_read),                                               //                          .read
		.av_readdata           (cpu_1_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_1_data_master_write),                                              //                          .write
		.av_writedata          (cpu_1_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_1_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_0_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ins_mem_0_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ins_mem_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ins_mem_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ins_mem_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ins_mem_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ins_mem_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ins_mem_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ins_mem_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atob_0_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                   //                    reset.reset
		.uav_address           (atob_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atob_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atob_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atob_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atob_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atob_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atob_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atob_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atob_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atob_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atob_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (atob_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (atob_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (atob_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atob_0_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                       //                    reset.reset
		.uav_address           (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (atob_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (atob_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (atob_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (atob_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (atob_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atob_0_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                    //                    reset.reset
		.uav_address           (atob_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atob_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atob_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atob_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atob_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atob_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atob_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atob_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atob_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atob_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atob_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (atob_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (atob_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (atob_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atob_1_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                   //                    reset.reset
		.uav_address           (atob_1_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atob_1_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atob_1_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atob_1_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atob_1_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atob_1_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atob_1_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atob_1_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atob_1_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atob_1_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atob_1_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (atob_1_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (atob_1_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (atob_1_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atob_1_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                       //                    reset.reset
		.uav_address           (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (atob_1_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (atob_1_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (atob_1_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (atob_1_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (atob_1_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atob_1_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                    //                    reset.reset
		.uav_address           (atob_1_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atob_1_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atob_1_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atob_1_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atob_1_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atob_1_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atob_1_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atob_1_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atob_1_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atob_1_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atob_1_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (atob_1_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (atob_1_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (atob_1_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atob_2_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                   //                    reset.reset
		.uav_address           (atob_2_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atob_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atob_2_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atob_2_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atob_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atob_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atob_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atob_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atob_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atob_2_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atob_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (atob_2_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (atob_2_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (atob_2_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atob_2_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                       //                    reset.reset
		.uav_address           (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (atob_2_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (atob_2_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (atob_2_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (atob_2_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (atob_2_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atob_2_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_007_reset_out_reset),                                    //                    reset.reset
		.uav_address           (atob_2_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atob_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atob_2_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atob_2_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atob_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atob_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atob_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atob_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atob_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atob_2_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atob_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (atob_2_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (atob_2_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (atob_2_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atod_0_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_013_reset_out_reset),                                   //                    reset.reset
		.uav_address           (atod_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atod_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atod_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atod_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atod_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atod_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atod_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atod_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atod_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atod_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atod_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (atod_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (atod_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (atod_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atod_0_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_013_reset_out_reset),                                    //                    reset.reset
		.uav_address           (atod_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atod_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atod_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atod_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atod_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atod_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atod_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atod_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atod_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atod_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atod_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (atod_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (atod_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (atod_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atod_0_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_013_reset_out_reset),                                       //                    reset.reset
		.uav_address           (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (atod_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (atod_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (atod_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (atod_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (atod_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atoe_0_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_014_reset_out_reset),                                   //                    reset.reset
		.uav_address           (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (atoe_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (atoe_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (atoe_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atoe_0_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_014_reset_out_reset),                                    //                    reset.reset
		.uav_address           (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (atoe_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (atoe_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (atoe_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atoe_0_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_014_reset_out_reset),                                       //                    reset.reset
		.uav_address           (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (atoe_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (atoe_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (atoe_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (atoe_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (atoe_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atof_0_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_012_reset_out_reset),                                   //                    reset.reset
		.uav_address           (atof_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atof_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atof_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atof_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atof_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atof_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atof_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atof_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atof_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atof_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atof_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (atof_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (atof_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (atof_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atof_0_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_012_reset_out_reset),                                       //                    reset.reset
		.uav_address           (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (atof_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (atof_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (atof_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (atof_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (atof_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) atof_0_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_012_reset_out_reset),                                    //                    reset.reset
		.uav_address           (atof_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (atof_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (atof_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (atof_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (atof_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (atof_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (atof_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (atof_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (atof_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (atof_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (atof_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (atof_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (atof_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (atof_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ins_mem_5_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                      //                    reset.reset
		.uav_address           (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ins_mem_5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ins_mem_5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ins_mem_5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ins_mem_5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ins_mem_5_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ins_mem_5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ins_mem_5_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_5_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_5_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) etof_0_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_011_reset_out_reset),                                   //                    reset.reset
		.uav_address           (etof_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (etof_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (etof_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (etof_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (etof_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (etof_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (etof_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (etof_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (etof_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (etof_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (etof_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (etof_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (etof_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (etof_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) etof_0_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_011_reset_out_reset),                                       //                    reset.reset
		.uav_address           (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (etof_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (etof_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (etof_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (etof_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (etof_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) etof_0_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_011_reset_out_reset),                                    //                    reset.reset
		.uav_address           (etof_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (etof_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (etof_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (etof_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (etof_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (etof_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (etof_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (etof_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (etof_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (etof_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (etof_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (etof_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (etof_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (etof_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_mem_5_s1_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                       //                    reset.reset
		.uav_address           (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_mem_5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (data_mem_5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (data_mem_5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (data_mem_5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (data_mem_5_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (data_mem_5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (data_mem_5_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_5_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_5_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_5_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_scale_timer_5_s1_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                               //                    reset.reset
		.uav_address           (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_scale_timer_5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_scale_timer_5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_scale_timer_5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_scale_timer_5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_scale_timer_5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                 //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_byteenable         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_mem_0_s1_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_mem_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (data_mem_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (data_mem_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (data_mem_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (data_mem_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (data_mem_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (data_mem_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_scale_timer_0_s1_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_scale_timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_scale_timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_scale_timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_scale_timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_scale_timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                 //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_byteenable         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ins_mem_4_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                      //                    reset.reset
		.uav_address           (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ins_mem_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ins_mem_4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ins_mem_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ins_mem_4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ins_mem_4_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ins_mem_4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ins_mem_4_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_4_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_4_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dtoe_0_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_010_reset_out_reset),                                   //                    reset.reset
		.uav_address           (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (dtoe_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (dtoe_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (dtoe_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dtoe_0_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_010_reset_out_reset),                                       //                    reset.reset
		.uav_address           (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (dtoe_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (dtoe_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (dtoe_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (dtoe_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (dtoe_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dtoe_0_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_010_reset_out_reset),                                    //                    reset.reset
		.uav_address           (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (dtoe_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (dtoe_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (dtoe_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_mem_4_s1_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                       //                    reset.reset
		.uav_address           (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_mem_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (data_mem_4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (data_mem_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (data_mem_4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (data_mem_4_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (data_mem_4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (data_mem_4_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_4_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_4_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_4_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_scale_timer_4_s1_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                               //                    reset.reset
		.uav_address           (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_scale_timer_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_scale_timer_4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_scale_timer_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_scale_timer_4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_scale_timer_4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                 //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_byteenable         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ins_mem_3_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                      //                    reset.reset
		.uav_address           (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ins_mem_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ins_mem_3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ins_mem_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ins_mem_3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ins_mem_3_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ins_mem_3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ins_mem_3_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_3_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_3_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ctod_0_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_009_reset_out_reset),                                   //                    reset.reset
		.uav_address           (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (ctod_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (ctod_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (ctod_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ctod_0_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_009_reset_out_reset),                                       //                    reset.reset
		.uav_address           (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ctod_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ctod_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ctod_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ctod_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ctod_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ctod_0_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_009_reset_out_reset),                                    //                    reset.reset
		.uav_address           (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (ctod_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (ctod_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (ctod_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_mem_3_s1_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                       //                    reset.reset
		.uav_address           (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_mem_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (data_mem_3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (data_mem_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (data_mem_3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (data_mem_3_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (data_mem_3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (data_mem_3_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_3_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_3_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_3_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_scale_timer_3_s1_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                               //                    reset.reset
		.uav_address           (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_scale_timer_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_scale_timer_3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_scale_timer_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_scale_timer_3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_scale_timer_3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                 //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_byteenable         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_mem_2_s1_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                       //                    reset.reset
		.uav_address           (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_mem_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (data_mem_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (data_mem_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (data_mem_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (data_mem_2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (data_mem_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (data_mem_2_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_2_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_2_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_2_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_scale_timer_2_s1_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                               //                    reset.reset
		.uav_address           (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_scale_timer_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_scale_timer_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_scale_timer_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_scale_timer_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_scale_timer_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                 //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_byteenable         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) btoc_0_in_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_008_reset_out_reset),                                   //                    reset.reset
		.uav_address           (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (btoc_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (btoc_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (btoc_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) btoc_0_out_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_008_reset_out_reset),                                    //                    reset.reset
		.uav_address           (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (btoc_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (btoc_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (btoc_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                      //              (terminated)
		.av_write              (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) btoc_0_in_csr_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_008_reset_out_reset),                                       //                    reset.reset
		.uav_address           (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (btoc_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (btoc_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (btoc_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (btoc_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (btoc_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ins_mem_2_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                      //                    reset.reset
		.uav_address           (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ins_mem_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ins_mem_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ins_mem_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ins_mem_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ins_mem_2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ins_mem_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ins_mem_2_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ins_mem_1_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address           (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ins_mem_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ins_mem_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ins_mem_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ins_mem_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ins_mem_1_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ins_mem_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ins_mem_1_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_1_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_mem_1_s1_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address           (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_mem_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (data_mem_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (data_mem_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (data_mem_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (data_mem_1_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (data_mem_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (data_mem_1_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_1_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_1_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (14),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_scale_timer_1_s1_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                               //                    reset.reset
		.uav_address           (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_scale_timer_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_scale_timer_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_scale_timer_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_scale_timer_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_scale_timer_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                 //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_byteenable         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                 //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                              //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                        //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                          //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                 //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_5_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_006_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (cpu_5_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_5_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_5_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_5_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_5_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_5_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_5_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_5_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_5_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_5_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_5_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_5_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_006_reset_out_reset),                                            // clk_reset.reset
		.av_address       (cpu_5_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_5_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_5_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_5_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_5_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_5_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_5_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_5_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_5_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_5_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_5_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_002_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_002_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_002_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_002_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_002_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_002_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_4_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_005_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (cpu_4_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_4_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_4_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_4_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_4_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_4_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_4_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_4_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_4_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_4_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_4_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_002_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_002_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_002_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_002_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_002_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_002_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_4_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_005_reset_out_reset),                                            // clk_reset.reset
		.av_address       (cpu_4_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_4_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_4_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_4_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_4_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_4_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_4_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_4_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_4_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_4_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_4_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_004_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_004_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_004_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_004_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_004_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_004_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (5),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_3_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_004_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (cpu_3_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_3_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_3_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_3_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_3_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_3_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_3_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_3_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_3_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_3_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_3_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_003_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_003_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_003_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_003_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_003_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_003_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (6),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_3_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_004_reset_out_reset),                                            // clk_reset.reset
		.av_address       (cpu_3_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_3_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_3_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_3_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_3_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_3_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_3_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_3_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_3_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_3_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_3_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_006_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_006_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_006_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_006_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_006_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_006_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (7),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_2_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                            // clk_reset.reset
		.av_address       (cpu_2_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_2_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_2_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_2_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_2_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_2_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_2_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_2_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_2_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_2_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_2_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_007_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_007_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_007_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_007_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_007_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_007_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (8),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_2_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (cpu_2_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_2_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_2_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_2_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_2_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_2_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_2_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_2_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_2_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_2_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_2_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_004_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_004_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_004_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_004_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_004_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_004_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (9),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_1_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_002_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (cpu_1_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_1_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_1_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_1_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_1_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_1_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_1_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_1_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_1_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_1_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_1_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_005_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_005_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_005_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_005_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_005_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_005_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (10),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_1_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.av_address       (cpu_1_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_1_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_1_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_1_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_1_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_1_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_1_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_1_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_1_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_1_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_1_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_010_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_010_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_010_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_010_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_010_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_010_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (11),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                       //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_011_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_011_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_011_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_011_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_011_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_011_src_ready)                                                     //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ins_mem_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                       //                .channel
		.rf_sink_ready           (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atob_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (atob_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atob_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atob_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atob_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atob_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atob_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atob_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atob_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atob_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atob_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atob_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atob_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atob_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atob_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atob_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atob_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                   //                .channel
		.rf_sink_ready           (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atob_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atob_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atob_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atob_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atob_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atob_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                             // clk_reset.reset
		.in_data           (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atob_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atob_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atob_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atob_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                       //                .channel
		.rf_sink_ready           (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atob_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (atob_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atob_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atob_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atob_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atob_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atob_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atob_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atob_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atob_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atob_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atob_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atob_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atob_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atob_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atob_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atob_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                    //                .channel
		.rf_sink_ready           (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atob_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atob_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atob_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atob_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atob_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atob_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                              // clk_reset.reset
		.in_data           (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atob_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atob_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atob_1_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (atob_1_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atob_1_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atob_1_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atob_1_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atob_1_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atob_1_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atob_1_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atob_1_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atob_1_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atob_1_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atob_1_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atob_1_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atob_1_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atob_1_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atob_1_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atob_1_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                   //                .channel
		.rf_sink_ready           (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atob_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atob_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atob_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atob_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atob_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atob_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                             // clk_reset.reset
		.in_data           (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atob_1_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atob_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atob_1_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atob_1_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_006_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_006_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_006_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_006_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_006_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_006_src_channel),                                                       //                .channel
		.rf_sink_ready           (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atob_1_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (atob_1_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atob_1_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atob_1_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atob_1_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atob_1_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atob_1_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atob_1_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atob_1_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atob_1_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atob_1_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atob_1_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atob_1_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atob_1_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atob_1_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atob_1_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atob_1_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_007_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_007_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_007_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_007_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_007_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_007_src_channel),                                                    //                .channel
		.rf_sink_ready           (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atob_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atob_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atob_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atob_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atob_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atob_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                              // clk_reset.reset
		.in_data           (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atob_1_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atob_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atob_2_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (atob_2_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atob_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atob_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atob_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atob_2_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atob_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atob_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atob_2_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atob_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atob_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atob_2_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atob_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atob_2_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atob_2_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atob_2_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atob_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                   //                .channel
		.rf_sink_ready           (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atob_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atob_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atob_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atob_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atob_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atob_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                             // clk_reset.reset
		.in_data           (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atob_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atob_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atob_2_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atob_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                       //                .channel
		.rf_sink_ready           (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atob_2_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_007_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (atob_2_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atob_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atob_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atob_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atob_2_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atob_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atob_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atob_2_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atob_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atob_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atob_2_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atob_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atob_2_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atob_2_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atob_2_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atob_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                    //                .channel
		.rf_sink_ready           (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atob_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atob_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atob_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atob_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atob_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atob_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_007_reset_out_reset),                                              // clk_reset.reset
		.in_data           (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atob_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atob_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atod_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_013_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (atod_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atod_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atod_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atod_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atod_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atod_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atod_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atod_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atod_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atod_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atod_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atod_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atod_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atod_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atod_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atod_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_011_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_011_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_011_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_011_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_011_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_011_src_channel),                                                   //                .channel
		.rf_sink_ready           (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_013_reset_out_reset),                                             // clk_reset.reset
		.in_data           (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atod_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atod_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_013_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (atod_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atod_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atod_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atod_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atod_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atod_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atod_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atod_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atod_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atod_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atod_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atod_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atod_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atod_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atod_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atod_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_012_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_012_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_012_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_012_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_012_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_012_src_channel),                                                    //                .channel
		.rf_sink_ready           (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_013_reset_out_reset),                                              // clk_reset.reset
		.in_data           (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atod_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atod_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_013_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_013_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_013_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_013_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_013_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_013_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_013_src_channel),                                                       //                .channel
		.rf_sink_ready           (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_013_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atoe_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_014_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atoe_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_014_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_014_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_014_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_014_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_014_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_014_src_channel),                                                   //                .channel
		.rf_sink_ready           (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_014_reset_out_reset),                                             // clk_reset.reset
		.in_data           (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atoe_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_014_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atoe_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_015_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_015_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_015_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_015_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_015_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_015_src_channel),                                                    //                .channel
		.rf_sink_ready           (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_014_reset_out_reset),                                              // clk_reset.reset
		.in_data           (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atoe_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_014_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_016_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_016_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_016_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_016_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_016_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_016_src_channel),                                                       //                .channel
		.rf_sink_ready           (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_014_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atof_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_012_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (atof_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atof_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atof_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atof_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atof_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atof_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atof_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atof_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atof_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atof_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atof_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atof_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atof_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atof_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atof_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atof_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_017_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_017_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_017_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_017_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_017_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_017_src_channel),                                                   //                .channel
		.rf_sink_ready           (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_012_reset_out_reset),                                             // clk_reset.reset
		.in_data           (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atof_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atof_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_012_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_018_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_018_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_018_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_018_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_018_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_018_src_channel),                                                       //                .channel
		.rf_sink_ready           (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_012_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) atof_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_012_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (atof_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (atof_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (atof_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (atof_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (atof_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (atof_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (atof_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (atof_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (atof_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (atof_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (atof_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (atof_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (atof_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (atof_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (atof_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (atof_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_019_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_019_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_019_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_019_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_019_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_019_src_channel),                                                    //                .channel
		.rf_sink_ready           (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (atof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (atof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (atof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (atof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (atof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (atof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_012_reset_out_reset),                                              // clk_reset.reset
		.in_data           (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (atof_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (atof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ins_mem_5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                   //                .channel
		.rf_sink_ready           (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_021_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_021_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_021_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_021_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_021_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_021_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) etof_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_011_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (etof_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (etof_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (etof_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (etof_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (etof_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (etof_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (etof_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (etof_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (etof_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (etof_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (etof_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (etof_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (etof_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (etof_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (etof_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (etof_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_022_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_022_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_022_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_022_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_022_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_022_src_channel),                                                   //                .channel
		.rf_sink_ready           (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (etof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (etof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (etof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (etof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (etof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (etof_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_011_reset_out_reset),                                             // clk_reset.reset
		.in_data           (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (etof_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (etof_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) etof_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_011_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (etof_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_023_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_023_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_023_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_023_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_023_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_023_src_channel),                                                       //                .channel
		.rf_sink_ready           (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_011_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) etof_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_011_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (etof_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (etof_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (etof_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (etof_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (etof_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (etof_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (etof_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (etof_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (etof_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (etof_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (etof_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (etof_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (etof_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (etof_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (etof_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (etof_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_024_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_024_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_024_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_024_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_024_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_024_src_channel),                                                    //                .channel
		.rf_sink_ready           (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (etof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (etof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (etof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (etof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (etof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (etof_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_011_reset_out_reset),                                              // clk_reset.reset
		.in_data           (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (etof_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (etof_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_mem_5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_mem_5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src7_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src7_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_002_src7_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src7_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src7_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src7_channel),                                                    //                .channel
		.rf_sink_ready           (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src8_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src8_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_002_src8_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src8_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src8_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src8_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src9_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src9_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src9_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src9_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src9_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src9_channel),                                                 //                .channel
		.rf_sink_ready           (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src10_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src10_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_002_src10_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src10_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src10_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src10_channel),                                                           //                .channel
		.rf_sink_ready           (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ins_mem_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src6_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src6_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_003_src6_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src6_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src6_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src6_channel),                                                   //                .channel
		.rf_sink_ready           (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_030_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_030_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_030_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_030_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_030_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_030_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dtoe_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_010_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dtoe_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_031_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_031_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_031_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_031_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_031_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_031_src_channel),                                                   //                .channel
		.rf_sink_ready           (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dtoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dtoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dtoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dtoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dtoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dtoe_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_010_reset_out_reset),                                             // clk_reset.reset
		.in_data           (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dtoe_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dtoe_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dtoe_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_010_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_032_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_032_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_032_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_032_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_032_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_032_src_channel),                                                       //                .channel
		.rf_sink_ready           (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_010_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dtoe_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_010_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dtoe_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_033_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_033_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_033_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_033_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_033_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_033_src_channel),                                                    //                .channel
		.rf_sink_ready           (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dtoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dtoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dtoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dtoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dtoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dtoe_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_010_reset_out_reset),                                              // clk_reset.reset
		.in_data           (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dtoe_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dtoe_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_mem_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_mem_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src10_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src10_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_004_src10_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src10_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src10_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src10_channel),                                                   //                .channel
		.rf_sink_ready           (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src11_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src11_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_004_src11_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src11_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src11_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src11_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src12_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src12_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_004_src12_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src12_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src12_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src12_channel),                                                //                .channel
		.rf_sink_ready           (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src13_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src13_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_004_src13_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src13_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src13_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src13_channel),                                                           //                .channel
		.rf_sink_ready           (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ins_mem_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src6_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src6_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_005_src6_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src6_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src6_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src6_channel),                                                   //                .channel
		.rf_sink_ready           (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_039_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_039_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_039_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_039_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_039_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_039_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ctod_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_009_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ctod_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_040_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_040_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_040_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_040_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_040_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_040_src_channel),                                                   //                .channel
		.rf_sink_ready           (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ctod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ctod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ctod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ctod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ctod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ctod_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_009_reset_out_reset),                                             // clk_reset.reset
		.in_data           (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ctod_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ctod_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ctod_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_009_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_041_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_041_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_041_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_041_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_041_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_041_src_channel),                                                       //                .channel
		.rf_sink_ready           (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_009_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ctod_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_009_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ctod_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_042_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_042_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_042_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_042_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_042_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_042_src_channel),                                                    //                .channel
		.rf_sink_ready           (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ctod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ctod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ctod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ctod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ctod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ctod_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_009_reset_out_reset),                                              // clk_reset.reset
		.in_data           (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ctod_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ctod_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_mem_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_mem_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src10_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src10_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_006_src10_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src10_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src10_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src10_channel),                                                   //                .channel
		.rf_sink_ready           (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src11_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src11_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_006_src11_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src11_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src11_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src11_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src12_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src12_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_006_src12_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src12_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src12_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src12_channel),                                                //                .channel
		.rf_sink_ready           (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_006_src13_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_006_src13_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_006_src13_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_006_src13_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_006_src13_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_006_src13_channel),                                                           //                .channel
		.rf_sink_ready           (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_mem_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src3_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src3_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_007_src3_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src3_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src3_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src3_channel),                                                    //                .channel
		.rf_sink_ready           (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_048_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_048_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_048_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_048_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_048_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_048_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src5_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src5_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_007_src5_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src5_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src5_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src5_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src6_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src6_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_007_src6_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src6_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src6_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src6_channel),                                                 //                .channel
		.rf_sink_ready           (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src7_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src7_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_007_src7_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src7_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src7_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src7_channel),                                                            //                .channel
		.rf_sink_ready           (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) btoc_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_008_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (btoc_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_052_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_052_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_052_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_052_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_052_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_052_src_channel),                                                   //                .channel
		.rf_sink_ready           (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (btoc_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (btoc_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (btoc_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (btoc_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (btoc_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (btoc_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_008_reset_out_reset),                                             // clk_reset.reset
		.in_data           (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (btoc_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (btoc_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) btoc_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_008_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (btoc_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_053_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_053_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_053_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_053_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_053_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_053_src_channel),                                                    //                .channel
		.rf_sink_ready           (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (btoc_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (btoc_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (btoc_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (btoc_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (btoc_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (btoc_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_008_reset_out_reset),                                              // clk_reset.reset
		.in_data           (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (btoc_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (btoc_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) btoc_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_008_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_054_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_054_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_054_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_054_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_054_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_054_src_channel),                                                       //                .channel
		.rf_sink_ready           (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_008_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ins_mem_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src7_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src7_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_008_src7_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src7_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src7_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src7_channel),                                                   //                .channel
		.rf_sink_ready           (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ins_mem_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_009_src12_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_009_src12_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_009_src12_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_009_src12_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_009_src12_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_009_src12_channel),                                                  //                .channel
		.rf_sink_ready           (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_057_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_057_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_057_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_057_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_057_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_057_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_mem_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_mem_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_010_src13_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_010_src13_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_010_src13_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_010_src13_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_010_src13_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_010_src13_channel),                                                   //                .channel
		.rf_sink_ready           (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_010_src14_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_010_src14_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_010_src14_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_010_src14_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_010_src14_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_010_src14_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_010_src15_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_010_src15_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_010_src15_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_010_src15_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_010_src15_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_010_src15_channel),                                                //                .channel
		.rf_sink_ready           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_010_src16_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_010_src16_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_010_src16_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_010_src16_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_010_src16_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_010_src16_channel),                                                           //                .channel
		.rf_sink_ready           (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_mem_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_mem_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_011_src19_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_011_src19_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_011_src19_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_011_src19_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_011_src19_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_011_src19_channel),                                                   //                .channel
		.rf_sink_ready           (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_011_src20_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_011_src20_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_011_src20_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_011_src20_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_011_src20_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_011_src20_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_011_src21_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_011_src21_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_011_src21_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_011_src21_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_011_src21_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_011_src21_channel),                                                //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (66),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_011_src22_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_011_src22_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_011_src22_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_011_src22_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_011_src22_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_011_src22_channel),                                                           //                .channel
		.rf_sink_ready           (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	SoC_addr_router addr_router (
		.sink_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	SoC_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_5_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_addr_router_002 addr_router_002 (
		.sink_ready         (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_5_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                     //          .valid
		.src_data           (addr_router_002_src_data),                                                      //          .data
		.src_channel        (addr_router_002_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_003 addr_router_003 (
		.sink_ready         (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_4_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                            //          .valid
		.src_data           (addr_router_003_src_data),                                                             //          .data
		.src_channel        (addr_router_003_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_addr_router_004 addr_router_004 (
		.sink_ready         (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_4_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                     //          .valid
		.src_data           (addr_router_004_src_data),                                                      //          .data
		.src_channel        (addr_router_004_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_005 addr_router_005 (
		.sink_ready         (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_3_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                            //          .valid
		.src_data           (addr_router_005_src_data),                                                             //          .data
		.src_channel        (addr_router_005_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_addr_router_006 addr_router_006 (
		.sink_ready         (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_3_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                     //          .valid
		.src_data           (addr_router_006_src_data),                                                      //          .data
		.src_channel        (addr_router_006_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_007 addr_router_007 (
		.sink_ready         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_007_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_007_src_valid),                                                     //          .valid
		.src_data           (addr_router_007_src_data),                                                      //          .data
		.src_channel        (addr_router_007_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_007_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_007_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_008 addr_router_008 (
		.sink_ready         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_008_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_008_src_valid),                                                            //          .valid
		.src_data           (addr_router_008_src_data),                                                             //          .data
		.src_channel        (addr_router_008_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_008_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_008_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_addr_router_009 addr_router_009 (
		.sink_ready         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_009_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_009_src_valid),                                                            //          .valid
		.src_data           (addr_router_009_src_data),                                                             //          .data
		.src_channel        (addr_router_009_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_009_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_009_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_addr_router_010 addr_router_010 (
		.sink_ready         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_010_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_010_src_valid),                                                     //          .valid
		.src_data           (addr_router_010_src_data),                                                      //          .data
		.src_channel        (addr_router_010_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_010_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_010_src_endofpacket)                                                //          .endofpacket
	);

	SoC_addr_router_011 addr_router_011 (
		.sink_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_011_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_011_src_valid),                                                     //          .valid
		.src_data           (addr_router_011_src_data),                                                      //          .data
		.src_channel        (addr_router_011_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_011_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_011_src_endofpacket)                                                //          .endofpacket
	);

	SoC_id_router id_router (
		.sink_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	SoC_id_router_001 id_router_001 (
		.sink_ready         (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ins_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                 //       src.ready
		.src_valid          (id_router_001_src_valid),                                                 //          .valid
		.src_data           (id_router_001_src_data),                                                  //          .data
		.src_channel        (id_router_001_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                            //          .endofpacket
	);

	SoC_id_router_002 id_router_002 (
		.sink_ready         (atob_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atob_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atob_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atob_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atob_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                              //       src.ready
		.src_valid          (id_router_002_src_valid),                                              //          .valid
		.src_data           (id_router_002_src_data),                                               //          .data
		.src_channel        (id_router_002_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_002 id_router_003 (
		.sink_ready         (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atob_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                  //       src.ready
		.src_valid          (id_router_003_src_valid),                                                  //          .valid
		.src_data           (id_router_003_src_data),                                                   //          .data
		.src_channel        (id_router_003_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_002 id_router_004 (
		.sink_ready         (atob_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atob_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atob_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atob_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atob_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                               //       src.ready
		.src_valid          (id_router_004_src_valid),                                               //          .valid
		.src_data           (id_router_004_src_data),                                                //          .data
		.src_channel        (id_router_004_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_002 id_router_005 (
		.sink_ready         (atob_1_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atob_1_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atob_1_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atob_1_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atob_1_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                              //       src.ready
		.src_valid          (id_router_005_src_valid),                                              //          .valid
		.src_data           (id_router_005_src_data),                                               //          .data
		.src_channel        (id_router_005_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_002 id_router_006 (
		.sink_ready         (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atob_1_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                  //       src.ready
		.src_valid          (id_router_006_src_valid),                                                  //          .valid
		.src_data           (id_router_006_src_data),                                                   //          .data
		.src_channel        (id_router_006_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_002 id_router_007 (
		.sink_ready         (atob_1_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atob_1_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atob_1_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atob_1_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atob_1_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                               //       src.ready
		.src_valid          (id_router_007_src_valid),                                               //          .valid
		.src_data           (id_router_007_src_data),                                                //          .data
		.src_channel        (id_router_007_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_002 id_router_008 (
		.sink_ready         (atob_2_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atob_2_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atob_2_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atob_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atob_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                              //       src.ready
		.src_valid          (id_router_008_src_valid),                                              //          .valid
		.src_data           (id_router_008_src_data),                                               //          .data
		.src_channel        (id_router_008_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_002 id_router_009 (
		.sink_ready         (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atob_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                  //       src.ready
		.src_valid          (id_router_009_src_valid),                                                  //          .valid
		.src_data           (id_router_009_src_data),                                                   //          .data
		.src_channel        (id_router_009_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_002 id_router_010 (
		.sink_ready         (atob_2_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atob_2_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atob_2_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atob_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atob_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                               //          .valid
		.src_data           (id_router_010_src_data),                                                //          .data
		.src_channel        (id_router_010_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_011 id_router_011 (
		.sink_ready         (atod_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atod_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atod_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atod_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atod_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                              //       src.ready
		.src_valid          (id_router_011_src_valid),                                              //          .valid
		.src_data           (id_router_011_src_data),                                               //          .data
		.src_channel        (id_router_011_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_011 id_router_012 (
		.sink_ready         (atod_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atod_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atod_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atod_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atod_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                               //       src.ready
		.src_valid          (id_router_012_src_valid),                                               //          .valid
		.src_data           (id_router_012_src_data),                                                //          .data
		.src_channel        (id_router_012_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_011 id_router_013 (
		.sink_ready         (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                  //       src.ready
		.src_valid          (id_router_013_src_valid),                                                  //          .valid
		.src_data           (id_router_013_src_data),                                                   //          .data
		.src_channel        (id_router_013_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_014 id_router_014 (
		.sink_ready         (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atoe_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                              //       src.ready
		.src_valid          (id_router_014_src_valid),                                              //          .valid
		.src_data           (id_router_014_src_data),                                               //          .data
		.src_channel        (id_router_014_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_014 id_router_015 (
		.sink_ready         (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atoe_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                               //       src.ready
		.src_valid          (id_router_015_src_valid),                                               //          .valid
		.src_data           (id_router_015_src_data),                                                //          .data
		.src_channel        (id_router_015_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_014 id_router_016 (
		.sink_ready         (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                  //       src.ready
		.src_valid          (id_router_016_src_valid),                                                  //          .valid
		.src_data           (id_router_016_src_data),                                                   //          .data
		.src_channel        (id_router_016_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_017 id_router_017 (
		.sink_ready         (atof_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atof_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atof_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atof_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atof_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                              //       src.ready
		.src_valid          (id_router_017_src_valid),                                              //          .valid
		.src_data           (id_router_017_src_data),                                               //          .data
		.src_channel        (id_router_017_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_017 id_router_018 (
		.sink_ready         (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                  //       src.ready
		.src_valid          (id_router_018_src_valid),                                                  //          .valid
		.src_data           (id_router_018_src_data),                                                   //          .data
		.src_channel        (id_router_018_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_017 id_router_019 (
		.sink_ready         (atof_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (atof_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (atof_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (atof_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (atof_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                               //       src.ready
		.src_valid          (id_router_019_src_valid),                                               //          .valid
		.src_data           (id_router_019_src_data),                                                //          .data
		.src_channel        (id_router_019_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_020 id_router_020 (
		.sink_ready         (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ins_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                 //       src.ready
		.src_valid          (id_router_020_src_valid),                                                 //          .valid
		.src_data           (id_router_020_src_data),                                                  //          .data
		.src_channel        (id_router_020_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                            //          .endofpacket
	);

	SoC_id_router_021 id_router_021 (
		.sink_ready         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_5_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                            //       src.ready
		.src_valid          (id_router_021_src_valid),                                                            //          .valid
		.src_data           (id_router_021_src_data),                                                             //          .data
		.src_channel        (id_router_021_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_022 id_router_022 (
		.sink_ready         (etof_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (etof_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (etof_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (etof_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (etof_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                              //       src.ready
		.src_valid          (id_router_022_src_valid),                                              //          .valid
		.src_data           (id_router_022_src_data),                                               //          .data
		.src_channel        (id_router_022_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_022 id_router_023 (
		.sink_ready         (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (etof_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                                  //       src.ready
		.src_valid          (id_router_023_src_valid),                                                  //          .valid
		.src_data           (id_router_023_src_data),                                                   //          .data
		.src_channel        (id_router_023_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_022 id_router_024 (
		.sink_ready         (etof_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (etof_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (etof_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (etof_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (etof_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                               //       src.ready
		.src_valid          (id_router_024_src_valid),                                               //          .valid
		.src_data           (id_router_024_src_data),                                                //          .data
		.src_channel        (id_router_024_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_025 id_router_025 (
		.sink_ready         (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_mem_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                  //       src.ready
		.src_valid          (id_router_025_src_valid),                                                  //          .valid
		.src_data           (id_router_025_src_data),                                                   //          .data
		.src_channel        (id_router_025_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_025 id_router_026 (
		.sink_ready         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_5_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_026_src_valid),                                                                  //          .valid
		.src_data           (id_router_026_src_data),                                                                   //          .data
		.src_channel        (id_router_026_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_025 id_router_027 (
		.sink_ready         (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                               //       src.ready
		.src_valid          (id_router_027_src_valid),                                               //          .valid
		.src_data           (id_router_027_src_data),                                                //          .data
		.src_channel        (id_router_027_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_025 id_router_028 (
		.sink_ready         (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_scale_timer_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                                          //       src.ready
		.src_valid          (id_router_028_src_valid),                                                          //          .valid
		.src_data           (id_router_028_src_data),                                                           //          .data
		.src_channel        (id_router_028_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                                     //          .endofpacket
	);

	SoC_id_router_029 id_router_029 (
		.sink_ready         (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ins_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                                 //       src.ready
		.src_valid          (id_router_029_src_valid),                                                 //          .valid
		.src_data           (id_router_029_src_data),                                                  //          .data
		.src_channel        (id_router_029_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                            //          .endofpacket
	);

	SoC_id_router_030 id_router_030 (
		.sink_ready         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_4_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                                            //       src.ready
		.src_valid          (id_router_030_src_valid),                                                            //          .valid
		.src_data           (id_router_030_src_data),                                                             //          .data
		.src_channel        (id_router_030_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_031 id_router_031 (
		.sink_ready         (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dtoe_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_031_src_ready),                                              //       src.ready
		.src_valid          (id_router_031_src_valid),                                              //          .valid
		.src_data           (id_router_031_src_data),                                               //          .data
		.src_channel        (id_router_031_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_031_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_031_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_031 id_router_032 (
		.sink_ready         (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dtoe_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_032_src_ready),                                                  //       src.ready
		.src_valid          (id_router_032_src_valid),                                                  //          .valid
		.src_data           (id_router_032_src_data),                                                   //          .data
		.src_channel        (id_router_032_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_032_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_032_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_031 id_router_033 (
		.sink_ready         (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dtoe_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_033_src_ready),                                               //       src.ready
		.src_valid          (id_router_033_src_valid),                                               //          .valid
		.src_data           (id_router_033_src_data),                                                //          .data
		.src_channel        (id_router_033_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_033_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_033_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_034 id_router_034 (
		.sink_ready         (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_mem_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_034_src_ready),                                                  //       src.ready
		.src_valid          (id_router_034_src_valid),                                                  //          .valid
		.src_data           (id_router_034_src_data),                                                   //          .data
		.src_channel        (id_router_034_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_034_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_034_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_034 id_router_035 (
		.sink_ready         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_4_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_035_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_035_src_valid),                                                                  //          .valid
		.src_data           (id_router_035_src_data),                                                                   //          .data
		.src_channel        (id_router_035_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_035_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_035_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_034 id_router_036 (
		.sink_ready         (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_036_src_ready),                                               //       src.ready
		.src_valid          (id_router_036_src_valid),                                               //          .valid
		.src_data           (id_router_036_src_data),                                                //          .data
		.src_channel        (id_router_036_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_036_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_036_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_034 id_router_037 (
		.sink_ready         (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_scale_timer_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_037_src_ready),                                                          //       src.ready
		.src_valid          (id_router_037_src_valid),                                                          //          .valid
		.src_data           (id_router_037_src_data),                                                           //          .data
		.src_channel        (id_router_037_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_037_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_037_src_endofpacket)                                                     //          .endofpacket
	);

	SoC_id_router_038 id_router_038 (
		.sink_ready         (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ins_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_038_src_ready),                                                 //       src.ready
		.src_valid          (id_router_038_src_valid),                                                 //          .valid
		.src_data           (id_router_038_src_data),                                                  //          .data
		.src_channel        (id_router_038_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_038_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_038_src_endofpacket)                                            //          .endofpacket
	);

	SoC_id_router_039 id_router_039 (
		.sink_ready         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_3_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_039_src_ready),                                                            //       src.ready
		.src_valid          (id_router_039_src_valid),                                                            //          .valid
		.src_data           (id_router_039_src_data),                                                             //          .data
		.src_channel        (id_router_039_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_039_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_039_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_040 id_router_040 (
		.sink_ready         (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ctod_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_040_src_ready),                                              //       src.ready
		.src_valid          (id_router_040_src_valid),                                              //          .valid
		.src_data           (id_router_040_src_data),                                               //          .data
		.src_channel        (id_router_040_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_040_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_040_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_040 id_router_041 (
		.sink_ready         (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ctod_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_041_src_ready),                                                  //       src.ready
		.src_valid          (id_router_041_src_valid),                                                  //          .valid
		.src_data           (id_router_041_src_data),                                                   //          .data
		.src_channel        (id_router_041_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_041_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_041_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_040 id_router_042 (
		.sink_ready         (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ctod_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_042_src_ready),                                               //       src.ready
		.src_valid          (id_router_042_src_valid),                                               //          .valid
		.src_data           (id_router_042_src_data),                                                //          .data
		.src_channel        (id_router_042_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_042_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_042_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_043 id_router_043 (
		.sink_ready         (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_mem_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_043_src_ready),                                                  //       src.ready
		.src_valid          (id_router_043_src_valid),                                                  //          .valid
		.src_data           (id_router_043_src_data),                                                   //          .data
		.src_channel        (id_router_043_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_043_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_043_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_043 id_router_044 (
		.sink_ready         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_3_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_044_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_044_src_valid),                                                                  //          .valid
		.src_data           (id_router_044_src_data),                                                                   //          .data
		.src_channel        (id_router_044_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_044_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_044_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_043 id_router_045 (
		.sink_ready         (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_045_src_ready),                                               //       src.ready
		.src_valid          (id_router_045_src_valid),                                               //          .valid
		.src_data           (id_router_045_src_data),                                                //          .data
		.src_channel        (id_router_045_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_045_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_045_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_043 id_router_046 (
		.sink_ready         (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_scale_timer_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_046_src_ready),                                                          //       src.ready
		.src_valid          (id_router_046_src_valid),                                                          //          .valid
		.src_data           (id_router_046_src_data),                                                           //          .data
		.src_channel        (id_router_046_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_046_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_046_src_endofpacket)                                                     //          .endofpacket
	);

	SoC_id_router_047 id_router_047 (
		.sink_ready         (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_047_src_ready),                                                  //       src.ready
		.src_valid          (id_router_047_src_valid),                                                  //          .valid
		.src_data           (id_router_047_src_data),                                                   //          .data
		.src_channel        (id_router_047_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_047_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_047_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_048 id_router_048 (
		.sink_ready         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_048_src_ready),                                                            //       src.ready
		.src_valid          (id_router_048_src_valid),                                                            //          .valid
		.src_data           (id_router_048_src_data),                                                             //          .data
		.src_channel        (id_router_048_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_048_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_048_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_047 id_router_049 (
		.sink_ready         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_049_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_049_src_valid),                                                                  //          .valid
		.src_data           (id_router_049_src_data),                                                                   //          .data
		.src_channel        (id_router_049_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_049_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_049_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_047 id_router_050 (
		.sink_ready         (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_050_src_ready),                                               //       src.ready
		.src_valid          (id_router_050_src_valid),                                               //          .valid
		.src_data           (id_router_050_src_data),                                                //          .data
		.src_channel        (id_router_050_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_050_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_050_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_047 id_router_051 (
		.sink_ready         (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_scale_timer_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_051_src_ready),                                                          //       src.ready
		.src_valid          (id_router_051_src_valid),                                                          //          .valid
		.src_data           (id_router_051_src_data),                                                           //          .data
		.src_channel        (id_router_051_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_051_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_051_src_endofpacket)                                                     //          .endofpacket
	);

	SoC_id_router_052 id_router_052 (
		.sink_ready         (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (btoc_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_052_src_ready),                                              //       src.ready
		.src_valid          (id_router_052_src_valid),                                              //          .valid
		.src_data           (id_router_052_src_data),                                               //          .data
		.src_channel        (id_router_052_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_052_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_052_src_endofpacket)                                         //          .endofpacket
	);

	SoC_id_router_052 id_router_053 (
		.sink_ready         (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (btoc_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_053_src_ready),                                               //       src.ready
		.src_valid          (id_router_053_src_valid),                                               //          .valid
		.src_data           (id_router_053_src_data),                                                //          .data
		.src_channel        (id_router_053_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_053_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_053_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_052 id_router_054 (
		.sink_ready         (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (btoc_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_054_src_ready),                                                  //       src.ready
		.src_valid          (id_router_054_src_valid),                                                  //          .valid
		.src_data           (id_router_054_src_data),                                                   //          .data
		.src_channel        (id_router_054_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_054_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_054_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_055 id_router_055 (
		.sink_ready         (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ins_mem_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_055_src_ready),                                                 //       src.ready
		.src_valid          (id_router_055_src_valid),                                                 //          .valid
		.src_data           (id_router_055_src_data),                                                  //          .data
		.src_channel        (id_router_055_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_055_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_055_src_endofpacket)                                            //          .endofpacket
	);

	SoC_id_router_056 id_router_056 (
		.sink_ready         (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ins_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_056_src_ready),                                                 //       src.ready
		.src_valid          (id_router_056_src_valid),                                                 //          .valid
		.src_data           (id_router_056_src_data),                                                  //          .data
		.src_channel        (id_router_056_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_056_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_056_src_endofpacket)                                            //          .endofpacket
	);

	SoC_id_router_057 id_router_057 (
		.sink_ready         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_057_src_ready),                                                            //       src.ready
		.src_valid          (id_router_057_src_valid),                                                            //          .valid
		.src_data           (id_router_057_src_data),                                                             //          .data
		.src_channel        (id_router_057_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_057_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_057_src_endofpacket)                                                       //          .endofpacket
	);

	SoC_id_router_058 id_router_058 (
		.sink_ready         (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_mem_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_058_src_ready),                                                  //       src.ready
		.src_valid          (id_router_058_src_valid),                                                  //          .valid
		.src_data           (id_router_058_src_data),                                                   //          .data
		.src_channel        (id_router_058_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_058_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_058_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_058 id_router_059 (
		.sink_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_059_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_059_src_valid),                                                                  //          .valid
		.src_data           (id_router_059_src_data),                                                                   //          .data
		.src_channel        (id_router_059_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_059_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_059_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_058 id_router_060 (
		.sink_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_060_src_ready),                                               //       src.ready
		.src_valid          (id_router_060_src_valid),                                               //          .valid
		.src_data           (id_router_060_src_data),                                                //          .data
		.src_channel        (id_router_060_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_060_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_060_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_058 id_router_061 (
		.sink_ready         (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_scale_timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_061_src_ready),                                                          //       src.ready
		.src_valid          (id_router_061_src_valid),                                                          //          .valid
		.src_data           (id_router_061_src_data),                                                           //          .data
		.src_channel        (id_router_061_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_061_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_061_src_endofpacket)                                                     //          .endofpacket
	);

	SoC_id_router_062 id_router_062 (
		.sink_ready         (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_mem_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_062_src_ready),                                                  //       src.ready
		.src_valid          (id_router_062_src_valid),                                                  //          .valid
		.src_data           (id_router_062_src_data),                                                   //          .data
		.src_channel        (id_router_062_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_062_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_062_src_endofpacket)                                             //          .endofpacket
	);

	SoC_id_router_062 id_router_063 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_063_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_063_src_valid),                                                                  //          .valid
		.src_data           (id_router_063_src_data),                                                                   //          .data
		.src_channel        (id_router_063_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_063_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_063_src_endofpacket)                                                             //          .endofpacket
	);

	SoC_id_router_062 id_router_064 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_064_src_ready),                                               //       src.ready
		.src_valid          (id_router_064_src_valid),                                               //          .valid
		.src_data           (id_router_064_src_data),                                                //          .data
		.src_channel        (id_router_064_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_064_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_064_src_endofpacket)                                          //          .endofpacket
	);

	SoC_id_router_062 id_router_065 (
		.sink_ready         (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_scale_timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_065_src_ready),                                                          //       src.ready
		.src_valid          (id_router_065_src_valid),                                                          //          .valid
		.src_data           (id_router_065_src_data),                                                           //          .data
		.src_channel        (id_router_065_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_065_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_065_src_endofpacket)                                                     //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.VALID_WIDTH               (66),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.VALID_WIDTH               (66),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_006_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.VALID_WIDTH               (66),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_005_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_003_src_data),           //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_003_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_003_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_003_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_003_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_003_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.VALID_WIDTH               (66),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_003 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_004_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_005_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_005_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_005_src_data),           //          .data
		.cmd_sink_channel       (addr_router_005_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_005_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_005_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_003_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_003_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_003_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_003_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_003_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_005_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_005_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_005_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_005_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_005_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_005_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_003_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_003_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_003_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_003_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_003_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_003_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_003_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.VALID_WIDTH               (66),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_004 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_008_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_008_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_008_src_data),           //          .data
		.cmd_sink_channel       (addr_router_008_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_008_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_008_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_004_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_004_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_004_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_004_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_004_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_008_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_008_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_008_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_008_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_008_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_008_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_004_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_004_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_004_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_004_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_004_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_004_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_004_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (66),
		.VALID_WIDTH               (66),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_005 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_002_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_009_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_009_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_009_src_data),           //          .data
		.cmd_sink_channel       (addr_router_009_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_009_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_009_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_005_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_005_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_005_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_005_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_005_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_009_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_009_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_009_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_009_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_009_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_009_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_005_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_005_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_005_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_005_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_005_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_005_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_005_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_1_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_004 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_3_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_005 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_4_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_006 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_5_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_006_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_007 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_1_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_007_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_008 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_2_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_1_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_008_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_009 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_3_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_2_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_009_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_010 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_3_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_4_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_010_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_011 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_4_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_5_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_011_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_012 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_5_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_0_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_012_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_013 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_3_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_013_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_014 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_4_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_014_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	SoC_cmd_xbar_demux cmd_xbar_demux (
		.clk                 (clk_clk),                            //        clk.clk
		.reset               (rst_controller_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_cmd_src_channel),            //           .channel
		.sink_data           (limiter_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_src18_endofpacket),   //           .endofpacket
		.src19_ready         (cmd_xbar_demux_src19_ready),         //      src19.ready
		.src19_valid         (cmd_xbar_demux_src19_valid),         //           .valid
		.src19_data          (cmd_xbar_demux_src19_data),          //           .data
		.src19_channel       (cmd_xbar_demux_src19_channel),       //           .channel
		.src19_startofpacket (cmd_xbar_demux_src19_startofpacket), //           .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_src19_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_006_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_006_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_002_src_ready),              //      sink.ready
		.sink_channel        (addr_router_002_src_channel),            //          .channel
		.sink_data           (addr_router_002_src_data),               //          .data
		.sink_startofpacket  (addr_router_002_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_002_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_002_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_002_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_002_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_002_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_002_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_002_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_002_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_002_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_002_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_002_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_002_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_002_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_002_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_002_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_002_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_002_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_002_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_002_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_002_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_002_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_002_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_002_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_002_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_002_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_002_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_002_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_002_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_002_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_002_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_002_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_002_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_002_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_002_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_002_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_002_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_002_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_002_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_002_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_002_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_002_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_002_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_002_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_002_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_002_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_002_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_002_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_002_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_002_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_002_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_002_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_002_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_002_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_002_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_002_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_002_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_002_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_002_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_002_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_002_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_002_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_002_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_002_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_002_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_002_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_002_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_002_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_002_src10_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                 (clk_clk),                                //        clk.clk
		.reset               (rst_controller_005_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_002_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_002_cmd_src_channel),            //           .channel
		.sink_data           (limiter_002_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_002_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_002_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_002_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_003_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_003_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_003_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_003_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_003_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_003_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_003_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_003_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_003_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_003_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_003_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_003_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_003_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_003_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_003_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_003_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_003_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_003_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_003_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_003_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_003_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_003_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_003_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_003_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_003_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_003_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_003_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_003_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_003_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_003_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_003_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_003_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_003_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_003_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_003_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_003_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_003_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_003_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_003_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_003_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_003_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_003_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_003_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_003_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_003_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_003_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_003_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_003_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_003_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_003_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_003_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_003_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_003_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_003_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_003_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_003_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_003_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_003_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_003_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_003_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_003_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_003_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_003_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_003_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_003_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_003_src10_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_005_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_004_src_ready),              //      sink.ready
		.sink_channel        (addr_router_004_src_channel),            //          .channel
		.sink_data           (addr_router_004_src_data),               //          .data
		.sink_startofpacket  (addr_router_004_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_004_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_004_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_004_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_004_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_004_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_004_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_004_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_004_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_004_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_004_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_004_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_004_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_004_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_004_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_004_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_004_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_004_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_004_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_004_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_004_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_004_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_004_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_004_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_004_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_004_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_004_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_004_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_004_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_004_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_004_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_004_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_004_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_004_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_004_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_004_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_004_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_004_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_004_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_004_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_004_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_004_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_004_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_004_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_004_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_004_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_004_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_004_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_004_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_004_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_004_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_004_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_004_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_004_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_004_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_004_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_004_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_004_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_004_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_004_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_004_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_004_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_004_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_004_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_004_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_004_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_004_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_004_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_004_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_004_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_004_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_004_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_004_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_004_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_004_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_004_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_004_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_004_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_004_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_004_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_004_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_004_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_004_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_004_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_004_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_004_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_004_src13_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_003 cmd_xbar_demux_005 (
		.clk                 (clk_clk),                                //        clk.clk
		.reset               (rst_controller_004_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_003_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_003_cmd_src_channel),            //           .channel
		.sink_data           (limiter_003_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_003_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_003_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_003_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_005_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_005_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_005_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_005_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_005_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_005_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_005_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_005_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_005_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_005_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_005_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_005_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_005_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_005_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_005_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_005_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_005_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_005_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_005_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_005_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_005_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_005_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_005_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_005_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_005_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_005_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_005_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_005_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_005_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_005_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_005_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_005_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_005_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_005_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_005_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_005_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_005_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_005_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_005_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_005_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_005_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_005_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_005_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_005_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_005_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_005_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_005_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_005_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_005_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_005_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_005_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_005_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_005_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_005_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_005_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_005_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_005_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_005_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_005_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_005_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_005_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_005_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_005_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_005_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_005_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_005_src10_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_004 cmd_xbar_demux_006 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_006_src_ready),              //      sink.ready
		.sink_channel        (addr_router_006_src_channel),            //          .channel
		.sink_data           (addr_router_006_src_data),               //          .data
		.sink_startofpacket  (addr_router_006_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_006_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_006_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_006_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_006_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_006_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_006_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_006_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_006_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_006_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_006_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_006_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_006_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_006_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_006_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_006_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_006_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_006_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_006_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_006_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_006_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_006_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_006_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_006_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_006_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_006_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_006_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_006_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_006_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_006_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_006_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_006_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_006_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_006_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_006_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_006_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_006_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_006_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_006_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_006_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_006_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_006_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_006_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_006_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_006_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_006_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_006_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_006_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_006_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_006_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_006_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_006_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_006_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_006_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_006_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_006_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_006_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_006_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_006_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_006_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_006_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_006_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_006_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_006_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_006_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_006_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_006_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_006_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_006_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_006_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_006_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_006_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_006_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_006_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_006_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_006_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_006_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_006_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_006_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_006_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_006_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_006_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_006_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_006_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_006_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_006_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_006_src13_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_002 cmd_xbar_demux_007 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_007_src_ready),              //      sink.ready
		.sink_channel        (addr_router_007_src_channel),            //          .channel
		.sink_data           (addr_router_007_src_data),               //          .data
		.sink_startofpacket  (addr_router_007_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_007_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_007_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_007_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_007_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_007_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_007_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_007_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_007_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_007_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_007_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_007_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_007_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_007_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_007_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_007_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_007_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_007_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_007_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_007_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_007_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_007_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_007_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_007_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_007_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_007_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_007_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_007_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_007_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_007_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_007_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_007_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_007_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_007_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_007_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_007_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_007_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_007_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_007_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_007_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_007_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_007_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_007_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_007_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_007_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_007_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_007_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_007_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_007_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_007_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_007_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_007_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_007_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_007_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_007_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_007_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_007_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_007_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_007_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_007_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_007_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_007_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_007_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_007_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_007_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_007_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_007_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_007_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_007_src10_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_001 cmd_xbar_demux_008 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_004_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_004_cmd_src_channel),           //           .channel
		.sink_data          (limiter_004_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_004_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_004_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_004_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_008_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_008_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_008_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_008_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_008_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_008_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_008_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_008_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_008_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_008_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_008_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_008_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_008_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_008_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_008_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_008_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_008_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_008_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_008_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_008_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_008_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_008_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_008_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_008_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_008_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_008_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_008_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_008_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_008_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_008_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_008_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_008_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_008_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_008_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_008_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_008_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_008_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_008_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_008_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_008_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_008_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_008_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_008_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_008_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_008_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_008_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_008_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_008_src7_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_009 cmd_xbar_demux_009 (
		.clk                 (clk_clk),                                //        clk.clk
		.reset               (rst_controller_002_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_005_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_005_cmd_src_channel),            //           .channel
		.sink_data           (limiter_005_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_005_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_005_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_005_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_009_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_009_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_009_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_009_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_009_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_009_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_009_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_009_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_009_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_009_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_009_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_009_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_009_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_009_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_009_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_009_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_009_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_009_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_009_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_009_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_009_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_009_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_009_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_009_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_009_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_009_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_009_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_009_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_009_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_009_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_009_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_009_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_009_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_009_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_009_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_009_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_009_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_009_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_009_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_009_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_009_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_009_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_009_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_009_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_009_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_009_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_009_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_009_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_009_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_009_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_009_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_009_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_009_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_009_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_009_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_009_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_009_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_009_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_009_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_009_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_009_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_009_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_009_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_009_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_009_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_009_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_009_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_009_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_009_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_009_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_009_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_009_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_009_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_009_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_009_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_009_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_009_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_009_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_009_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_009_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_009_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_009_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_009_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_009_src13_endofpacket)    //           .endofpacket
	);

	SoC_cmd_xbar_demux_010 cmd_xbar_demux_010 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_010_src_ready),              //      sink.ready
		.sink_channel        (addr_router_010_src_channel),            //          .channel
		.sink_data           (addr_router_010_src_data),               //          .data
		.sink_startofpacket  (addr_router_010_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_010_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_010_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_010_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_010_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_010_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_010_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_010_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_010_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_010_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_010_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_010_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_010_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_010_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_010_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_010_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_010_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_010_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_010_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_010_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_010_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_010_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_010_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_010_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_010_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_010_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_010_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_010_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_010_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_010_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_010_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_010_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_010_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_010_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_010_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_010_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_010_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_010_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_010_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_010_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_010_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_010_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_010_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_010_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_010_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_010_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_010_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_010_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_010_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_010_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_010_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_010_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_010_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_010_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_010_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_010_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_010_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_010_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_010_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_010_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_010_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_010_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_010_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_010_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_010_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_010_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_010_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_010_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_010_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_010_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_010_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_010_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_010_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_010_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_010_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_010_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_010_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_010_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_010_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_010_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_010_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_010_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_010_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_010_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_010_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_010_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_010_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_010_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_010_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_010_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_010_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_010_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_010_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_010_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_010_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_010_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_010_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_010_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_010_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_010_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_010_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_010_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_010_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_010_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_010_src16_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_demux_011 cmd_xbar_demux_011 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_011_src_ready),              //      sink.ready
		.sink_channel        (addr_router_011_src_channel),            //          .channel
		.sink_data           (addr_router_011_src_data),               //          .data
		.sink_startofpacket  (addr_router_011_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_011_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_011_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_011_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_011_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_011_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_011_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_011_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_011_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_011_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_011_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_011_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_011_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_011_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_011_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_011_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_011_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_011_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_011_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_011_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_011_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_011_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_011_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_011_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_011_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_011_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_011_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_011_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_011_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_011_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_011_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_011_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_011_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_011_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_011_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_011_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_011_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_011_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_011_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_011_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_011_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_011_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_011_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_011_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_011_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_011_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_011_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_011_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_011_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_011_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_011_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_011_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_011_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_011_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_011_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_011_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_011_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_011_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_011_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_011_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_011_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_011_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_011_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_011_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_011_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_011_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_011_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_011_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_011_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_011_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_011_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_011_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_011_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_011_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_011_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_011_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_011_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_011_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_011_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_011_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_011_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_011_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_011_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_011_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_011_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_011_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_011_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_011_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_011_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_011_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_011_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_011_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_011_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_011_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_011_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_011_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_011_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_011_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_011_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_011_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_011_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_011_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_011_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_011_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_011_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_011_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_011_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_011_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_011_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_011_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_011_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_011_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_011_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_011_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_011_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_011_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_011_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_011_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_011_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_011_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_011_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_011_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_011_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_011_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_011_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_011_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_011_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_011_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_011_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_011_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_011_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_011_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_011_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_011_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_011_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_011_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_011_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_011_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_011_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_011_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_011_src22_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_011_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_011_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_011_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_011_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_010_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_010_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_010_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_010_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src1_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src1_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src1_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src1_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src1_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_010_src1_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_010_src1_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_010_src1_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_010_src1_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src2_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src2_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src2_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src2_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src2_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src2_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_004 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src2_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_010_src2_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_010_src2_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_010_src2_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_010_src2_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_010_src2_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src3_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src3_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src3_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src3_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src3_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src3_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_005 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src3_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_010_src3_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_010_src3_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_010_src3_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_010_src3_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_010_src3_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_010_src3_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src4_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src4_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src4_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src4_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src4_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src4_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_006 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src4_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_010_src4_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_010_src4_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_010_src4_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_010_src4_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_010_src4_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_010_src4_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src5_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src5_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src5_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src5_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src5_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src5_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_007 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src7_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src7_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src7_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src7_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src7_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src7_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src5_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_010_src5_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_010_src5_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_010_src5_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_010_src5_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_010_src5_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_010_src5_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src6_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src6_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src6_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src6_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src6_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src6_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_008 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src8_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src8_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src8_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src8_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src8_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src8_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src6_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src6_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src6_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src6_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src6_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src6_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_010_src6_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_010_src6_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_010_src6_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_010_src6_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_010_src6_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_010_src6_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src7_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src7_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src7_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src7_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src7_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src7_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_009 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src9_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src9_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src9_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src9_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src9_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src9_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src7_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src7_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src7_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src7_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src7_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src7_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_010_src7_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_010_src7_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_010_src7_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_010_src7_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_010_src7_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_010_src7_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src8_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src8_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src8_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src8_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src8_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src8_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_010 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src10_ready),            //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src10_valid),            //          .valid
		.sink0_channel       (cmd_xbar_demux_src10_channel),          //          .channel
		.sink0_data          (cmd_xbar_demux_src10_data),             //          .data
		.sink0_startofpacket (cmd_xbar_demux_src10_startofpacket),    //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src10_endofpacket),      //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_009_src8_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_009_src8_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_009_src8_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_009_src8_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_009_src8_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_009_src8_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_010_src8_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_010_src8_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_010_src8_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_010_src8_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_010_src8_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_010_src8_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src9_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src9_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src9_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src9_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src9_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src9_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_011 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_013_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_011_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_011_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_011_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_011_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_011_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_011_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src11_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src11_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src11_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src11_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src11_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src11_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_005_src0_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_005_src0_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_005_src0_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_005_src0_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_005_src0_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_005_src0_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_006_src0_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_006_src0_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_006_src0_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_006_src0_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_006_src0_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_006_src0_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src10_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src10_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src10_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src10_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src10_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src10_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_012 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_013_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_012_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_012_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_012_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_012_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_012_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_012_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src12_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src12_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src12_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src12_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src12_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src12_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_005_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_005_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_005_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_005_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_005_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_005_src1_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_006_src1_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_006_src1_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_006_src1_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_006_src1_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_006_src1_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_006_src1_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src11_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src11_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src11_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src11_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src11_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src11_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_013 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_013_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_013_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_013_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_013_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_013_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_013_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_013_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src13_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src13_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src13_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src13_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src13_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src13_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_005_src2_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_005_src2_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_005_src2_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_005_src2_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_005_src2_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_005_src2_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_006_src2_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_006_src2_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_006_src2_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_006_src2_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_006_src2_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_006_src2_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src12_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src12_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src12_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src12_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src12_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src12_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_014 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_014_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_014_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_014_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_014_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_014_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_014_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_014_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src14_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src14_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src14_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src14_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src14_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src14_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src0_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src0_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src0_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_003_src0_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src0_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src0_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src0_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src0_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_004_src0_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src0_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src13_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src13_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src13_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src13_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src13_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src13_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_015 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_014_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_015_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_015_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_015_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_015_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_015_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_015_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src15_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src15_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src15_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src15_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src15_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src15_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_003_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src1_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src1_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src1_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_004_src1_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src1_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src1_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src14_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src14_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src14_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src14_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src14_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src14_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_016 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_014_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_016_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_016_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_016_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_016_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_016_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_016_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src16_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src16_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src16_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src16_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src16_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src16_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src2_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src2_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src2_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_003_src2_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src2_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src2_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src2_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src2_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src2_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_004_src2_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src2_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src2_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src15_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src15_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src15_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src15_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src15_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src15_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_017 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_012_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_017_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_017_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_017_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_017_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_017_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_017_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src17_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src17_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src17_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src17_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src17_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src17_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src0_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src0_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src0_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_002_src0_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src0_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src16_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src16_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src16_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src16_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src16_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src16_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_018 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_012_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_018_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_018_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_018_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_018_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_018_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_018_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src18_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src18_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src18_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src18_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src18_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src18_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src1_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src1_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src1_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_002_src1_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src1_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src17_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src17_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src17_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src17_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src17_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src17_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_019 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_012_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_019_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_019_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_019_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_019_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_019_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_019_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src19_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src19_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src19_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src19_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src19_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src19_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src2_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src2_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src2_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_002_src2_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src2_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_011_src18_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_011_src18_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_011_src18_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_011_src18_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_011_src18_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_011_src18_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_021 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_021_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_021_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_021_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_021_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_021_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_021_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src4_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src3_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_022 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_011_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_022_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_022_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_022_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_022_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_022_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_022_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src5_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src4_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src3_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src3_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src3_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src3_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src3_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src3_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src3_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src3_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_004_src3_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src3_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src3_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_023 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_011_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_023_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_023_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_023_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_023_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_023_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_023_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src6_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src5_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src4_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src4_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src4_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src4_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src4_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src4_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src4_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src4_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src4_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_004_src4_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src4_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src4_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_024 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_011_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_024_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_024_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_024_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_024_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_024_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_024_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src7_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src6_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src6_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src6_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src6_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src6_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src6_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src5_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src5_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src5_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src5_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src5_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src5_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src5_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src5_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src5_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_004_src5_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src5_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src5_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_030 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_030_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_030_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_030_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_030_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_030_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_030_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src7_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src7_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src7_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src7_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src7_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src7_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_004_src6_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_004_src6_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_004_src6_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_004_src6_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_004_src6_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_004_src6_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_031 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_010_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_031_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_031_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_031_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_031_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_031_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_031_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src8_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src8_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src8_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src8_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src8_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src8_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_004_src7_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_004_src7_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_004_src7_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_004_src7_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_004_src7_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_004_src7_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_005_src3_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_005_src3_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_005_src3_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_005_src3_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_005_src3_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_005_src3_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_006_src3_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_006_src3_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_006_src3_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_006_src3_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_006_src3_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_006_src3_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_032 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_010_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_032_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_032_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_032_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_032_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_032_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_032_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src9_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src9_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src9_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src9_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src9_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src9_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_004_src8_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_004_src8_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_004_src8_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_004_src8_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_004_src8_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_004_src8_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_005_src4_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_005_src4_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_005_src4_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_005_src4_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_005_src4_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_005_src4_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_006_src4_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_006_src4_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_006_src4_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_006_src4_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_006_src4_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_006_src4_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_033 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_010_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_033_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_033_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_033_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_033_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_033_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_033_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src10_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src10_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src10_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src10_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src10_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src10_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_004_src9_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_004_src9_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_004_src9_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_004_src9_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_004_src9_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_004_src9_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_005_src5_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_005_src5_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_005_src5_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_005_src5_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_005_src5_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_005_src5_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_006_src5_ready),          //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_006_src5_valid),          //          .valid
		.sink3_channel       (cmd_xbar_demux_006_src5_channel),        //          .channel
		.sink3_data          (cmd_xbar_demux_006_src5_data),           //          .data
		.sink3_startofpacket (cmd_xbar_demux_006_src5_startofpacket),  //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_006_src5_endofpacket)     //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_039 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_039_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_039_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_039_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_039_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_039_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_039_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_005_src7_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_005_src7_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_005_src7_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_005_src7_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_005_src7_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_005_src7_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_006_src6_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_006_src6_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_006_src6_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_006_src6_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_006_src6_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_006_src6_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_040 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_009_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_040_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_040_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_040_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_040_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_040_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_040_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_005_src8_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_005_src8_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_005_src8_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_005_src8_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_005_src8_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_005_src8_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_006_src7_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_006_src7_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_006_src7_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_006_src7_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_006_src7_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_006_src7_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_007_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_007_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_007_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_007_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_008_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_008_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_008_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_008_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_041 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_009_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_041_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_041_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_041_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_041_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_041_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_041_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_005_src9_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_005_src9_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_005_src9_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_005_src9_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_005_src9_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_005_src9_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_006_src8_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_006_src8_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_006_src8_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_006_src8_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_006_src8_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_006_src8_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_007_src1_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_007_src1_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_007_src1_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_007_src1_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_008_src1_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_008_src1_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_008_src1_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_008_src1_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_042 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_009_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_042_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_042_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_042_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_042_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_042_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_042_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_005_src10_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_005_src10_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_005_src10_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_005_src10_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_005_src10_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_005_src10_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_006_src9_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_006_src9_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_006_src9_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_006_src9_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_006_src9_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_006_src9_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_007_src2_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_007_src2_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_007_src2_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_007_src2_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_007_src2_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_007_src2_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_008_src2_ready),          //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_008_src2_valid),          //          .valid
		.sink3_channel       (cmd_xbar_demux_008_src2_channel),        //          .channel
		.sink3_data          (cmd_xbar_demux_008_src2_data),           //          .data
		.sink3_startofpacket (cmd_xbar_demux_008_src2_startofpacket),  //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_008_src2_endofpacket)     //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_048 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_048_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_048_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_048_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_048_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_048_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_048_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_007_src4_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_007_src4_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_007_src4_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_007_src4_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_007_src4_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_007_src4_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_008_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_008_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_008_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_008_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_008_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_008_src3_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_052 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_008_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_052_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_052_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_052_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_052_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_052_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_052_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_007_src8_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_007_src8_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_007_src8_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_007_src8_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_007_src8_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_007_src8_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_008_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_008_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_008_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_008_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_008_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_008_src4_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_009_src9_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_009_src9_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_009_src9_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_009_src9_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_009_src9_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_009_src9_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_010_src9_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_010_src9_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_010_src9_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_010_src9_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_010_src9_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_010_src9_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_053 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_008_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_053_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_053_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_053_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_053_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_053_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_053_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_007_src9_ready),          //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_007_src9_valid),          //          .valid
		.sink0_channel       (cmd_xbar_demux_007_src9_channel),        //          .channel
		.sink0_data          (cmd_xbar_demux_007_src9_data),           //          .data
		.sink0_startofpacket (cmd_xbar_demux_007_src9_startofpacket),  //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_007_src9_endofpacket),    //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_008_src5_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_008_src5_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_008_src5_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_008_src5_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_008_src5_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_008_src5_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_009_src10_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_009_src10_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_009_src10_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_009_src10_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_009_src10_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_009_src10_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_010_src10_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_010_src10_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_010_src10_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_010_src10_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_010_src10_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_010_src10_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux_002 cmd_xbar_mux_054 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_008_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_054_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_054_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_054_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_054_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_054_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_054_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_007_src10_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_007_src10_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_007_src10_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_007_src10_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_007_src10_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_007_src10_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_008_src6_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_008_src6_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_008_src6_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_008_src6_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_008_src6_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_008_src6_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_009_src11_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_009_src11_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_009_src11_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_009_src11_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_009_src11_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_009_src11_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_010_src11_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_010_src11_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_010_src11_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_010_src11_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_010_src11_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_010_src11_endofpacket)    //          .endofpacket
	);

	SoC_cmd_xbar_mux cmd_xbar_mux_057 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_057_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_057_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_057_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_057_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_057_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_057_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_009_src13_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_009_src13_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_009_src13_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_009_src13_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_009_src13_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_009_src13_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_010_src12_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_010_src12_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_010_src12_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_010_src12_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_010_src12_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_010_src12_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_002_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_003_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_003_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_003_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_003_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_003_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_003_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_004_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_004_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_004_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_004_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_004_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_004_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_004_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_004_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_004_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_004_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_004_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_004_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_005_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_005_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_005_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_005_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_005_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_005_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_005_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_005_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_005_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_005_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_005_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_005_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_006_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_006_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_006_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_006_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_006_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_006_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_006_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_006_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_006_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_006_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_006_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_006_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_007_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_007_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_007_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_007_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_007_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_007_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_007_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_007_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_007_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_007_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_007_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_007_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_008_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_008_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_008_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_008_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_008_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_008_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_008_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_008_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_008_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_008_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_008_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_008_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_009_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_009_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_009_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_009_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_009_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_009_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_009_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_009_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_009_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_009_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_009_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_009_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_007_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_010_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_010_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_010_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_010_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_010_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_010_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_010_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_010_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_010_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_010_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_010_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_011_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_011_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_011_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_011_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_011_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_011_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_011_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_011_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_011_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_011_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_011_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_011_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_011_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_011_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_011_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_011_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_011_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_012_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_012_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_012_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_012_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_012_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_012_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_012_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_012_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_012_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_012_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_012_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_012_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_012_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_012_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_013_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_013_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_013_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_013_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_013_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_013_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_013_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_013_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_013_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_013_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_013_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_013_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_013_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_013_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_013_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_014 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_014_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_014_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_014_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_014_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_014_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_014_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_014_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_014_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_014_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_014_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_014_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_014_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_014_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_014_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_014_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_014_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_014_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_015 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_015_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_015_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_015_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_015_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_015_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_015_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_015_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_015_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_015_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_015_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_015_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_015_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_015_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_015_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_016 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_014_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_016_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_016_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_016_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_016_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_016_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_016_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_016_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_016_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_016_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_016_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_016_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_016_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_016_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_016_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_016_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_016_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_016_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_016_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_017 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_017_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_017_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_017_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_017_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_017_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_017_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_017_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_017_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_017_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_017_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_017_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_017_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_017_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_017_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_017_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_017_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_017_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_017_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_018 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_018_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_018_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_018_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_018_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_018_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_018_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_018_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_018_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_018_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_018_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_018_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_018_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_018_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_018_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_018_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_018_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_018_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_018_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_019 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_012_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_019_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_019_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_019_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_019_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_019_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_019_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_019_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_019_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_019_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_019_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_019_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_019_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_019_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_019_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_019_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_019_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_019_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_019_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_020 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_021 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_021_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_021_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_021_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_021_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_021_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_021_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_022 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_022_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_022_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_022_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_022_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_022_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_022_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_022_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_022_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_022_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_022_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_022_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_022_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_022_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_022_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_022_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_022_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_022_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_022_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_023 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_023_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_023_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_023_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_023_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_023_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_023_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_023_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_023_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_023_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_023_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_023_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_023_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_023_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_023_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_023_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_023_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_023_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_023_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_024 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_011_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_024_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_024_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_024_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_024_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_024_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_024_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_024_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_024_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_024_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_024_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_024_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_024_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_024_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_024_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_024_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_024_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_024_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_024_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_025 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_026 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_027 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_028 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_029 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_029_src_ready),               //      sink.ready
		.sink_channel       (id_router_029_src_channel),             //          .channel
		.sink_data          (id_router_029_src_data),                //          .data
		.sink_startofpacket (id_router_029_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_029_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_029_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_030 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_030_src_ready),               //      sink.ready
		.sink_channel       (id_router_030_src_channel),             //          .channel
		.sink_data          (id_router_030_src_data),                //          .data
		.sink_startofpacket (id_router_030_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_030_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_030_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_030_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_030_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_030_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_030_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_030_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_030_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_031 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_031_src_ready),               //      sink.ready
		.sink_channel       (id_router_031_src_channel),             //          .channel
		.sink_data          (id_router_031_src_data),                //          .data
		.sink_startofpacket (id_router_031_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_031_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_031_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_031_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_031_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_031_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_031_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_031_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_031_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_031_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_031_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_031_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_031_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_031_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_031_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_031_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_031_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_031_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_031_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_031_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_031_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_031_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_032 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_032_src_ready),               //      sink.ready
		.sink_channel       (id_router_032_src_channel),             //          .channel
		.sink_data          (id_router_032_src_data),                //          .data
		.sink_startofpacket (id_router_032_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_032_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_032_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_032_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_032_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_032_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_032_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_032_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_032_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_032_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_032_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_032_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_032_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_032_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_032_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_032_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_032_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_032_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_032_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_032_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_032_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_032_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_032_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_033 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_010_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_033_src_ready),               //      sink.ready
		.sink_channel       (id_router_033_src_channel),             //          .channel
		.sink_data          (id_router_033_src_data),                //          .data
		.sink_startofpacket (id_router_033_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_033_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_033_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_033_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_033_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_033_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_033_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_033_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_033_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_033_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_033_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_033_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_033_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_033_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_033_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_033_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_033_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_033_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_033_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_033_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_033_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_033_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_033_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_034 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_034_src_ready),               //      sink.ready
		.sink_channel       (id_router_034_src_channel),             //          .channel
		.sink_data          (id_router_034_src_data),                //          .data
		.sink_startofpacket (id_router_034_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_034_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_034_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_034_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_034_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_035 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_035_src_ready),               //      sink.ready
		.sink_channel       (id_router_035_src_channel),             //          .channel
		.sink_data          (id_router_035_src_data),                //          .data
		.sink_startofpacket (id_router_035_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_035_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_035_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_035_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_035_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_036 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_036_src_ready),               //      sink.ready
		.sink_channel       (id_router_036_src_channel),             //          .channel
		.sink_data          (id_router_036_src_data),                //          .data
		.sink_startofpacket (id_router_036_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_036_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_036_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_036_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_037 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_037_src_ready),               //      sink.ready
		.sink_channel       (id_router_037_src_channel),             //          .channel
		.sink_data          (id_router_037_src_data),                //          .data
		.sink_startofpacket (id_router_037_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_037_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_037_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_037_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_037_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_038 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_038_src_ready),               //      sink.ready
		.sink_channel       (id_router_038_src_channel),             //          .channel
		.sink_data          (id_router_038_src_data),                //          .data
		.sink_startofpacket (id_router_038_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_038_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_038_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_038_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_038_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_038_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_038_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_038_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_039 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_039_src_ready),               //      sink.ready
		.sink_channel       (id_router_039_src_channel),             //          .channel
		.sink_data          (id_router_039_src_data),                //          .data
		.sink_startofpacket (id_router_039_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_039_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_039_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_039_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_039_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_039_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_039_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_039_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_039_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_039_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_039_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_039_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_039_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_039_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_040 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_040_src_ready),               //      sink.ready
		.sink_channel       (id_router_040_src_channel),             //          .channel
		.sink_data          (id_router_040_src_data),                //          .data
		.sink_startofpacket (id_router_040_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_040_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_040_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_040_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_040_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_040_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_040_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_040_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_040_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_040_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_040_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_040_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_040_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_040_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_040_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_040_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_040_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_040_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_040_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_040_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_040_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_040_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_040_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_040_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_040_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_040_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_041 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_041_src_ready),               //      sink.ready
		.sink_channel       (id_router_041_src_channel),             //          .channel
		.sink_data          (id_router_041_src_data),                //          .data
		.sink_startofpacket (id_router_041_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_041_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_041_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_041_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_041_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_041_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_041_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_041_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_041_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_041_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_041_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_041_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_041_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_041_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_041_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_041_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_041_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_041_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_041_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_041_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_041_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_041_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_041_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_041_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_041_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_041_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_042 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_009_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_042_src_ready),               //      sink.ready
		.sink_channel       (id_router_042_src_channel),             //          .channel
		.sink_data          (id_router_042_src_data),                //          .data
		.sink_startofpacket (id_router_042_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_042_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_042_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_042_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_042_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_042_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_042_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_042_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_042_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_042_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_042_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_042_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_042_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_042_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_042_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_042_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_042_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_042_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_042_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_042_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_042_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_042_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_042_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_043 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_043_src_ready),               //      sink.ready
		.sink_channel       (id_router_043_src_channel),             //          .channel
		.sink_data          (id_router_043_src_data),                //          .data
		.sink_startofpacket (id_router_043_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_043_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_043_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_043_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_043_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_044 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_044_src_ready),               //      sink.ready
		.sink_channel       (id_router_044_src_channel),             //          .channel
		.sink_data          (id_router_044_src_data),                //          .data
		.sink_startofpacket (id_router_044_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_044_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_044_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_044_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_044_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_045 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_045_src_ready),               //      sink.ready
		.sink_channel       (id_router_045_src_channel),             //          .channel
		.sink_data          (id_router_045_src_data),                //          .data
		.sink_startofpacket (id_router_045_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_045_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_045_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_045_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_045_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_046 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_046_src_ready),               //      sink.ready
		.sink_channel       (id_router_046_src_channel),             //          .channel
		.sink_data          (id_router_046_src_data),                //          .data
		.sink_startofpacket (id_router_046_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_046_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_046_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_046_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_046_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_047 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_047_src_ready),               //      sink.ready
		.sink_channel       (id_router_047_src_channel),             //          .channel
		.sink_data          (id_router_047_src_data),                //          .data
		.sink_startofpacket (id_router_047_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_047_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_047_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_047_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_047_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_047_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_047_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_047_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_048 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_048_src_ready),               //      sink.ready
		.sink_channel       (id_router_048_src_channel),             //          .channel
		.sink_data          (id_router_048_src_data),                //          .data
		.sink_startofpacket (id_router_048_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_048_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_048_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_048_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_048_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_048_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_048_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_048_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_048_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_048_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_048_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_048_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_048_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_048_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_049 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_049_src_ready),               //      sink.ready
		.sink_channel       (id_router_049_src_channel),             //          .channel
		.sink_data          (id_router_049_src_data),                //          .data
		.sink_startofpacket (id_router_049_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_049_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_049_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_049_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_049_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_049_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_049_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_049_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_050 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_050_src_ready),               //      sink.ready
		.sink_channel       (id_router_050_src_channel),             //          .channel
		.sink_data          (id_router_050_src_data),                //          .data
		.sink_startofpacket (id_router_050_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_050_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_050_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_050_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_050_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_050_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_050_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_050_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_051 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_051_src_ready),               //      sink.ready
		.sink_channel       (id_router_051_src_channel),             //          .channel
		.sink_data          (id_router_051_src_data),                //          .data
		.sink_startofpacket (id_router_051_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_051_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_051_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_051_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_051_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_051_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_051_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_051_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_052 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_052_src_ready),               //      sink.ready
		.sink_channel       (id_router_052_src_channel),             //          .channel
		.sink_data          (id_router_052_src_data),                //          .data
		.sink_startofpacket (id_router_052_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_052_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_052_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_052_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_052_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_052_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_052_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_052_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_052_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_052_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_052_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_052_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_052_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_052_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_052_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_052_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_052_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_052_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_052_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_052_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_052_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_052_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_052_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_052_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_052_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_052_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_053 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_053_src_ready),               //      sink.ready
		.sink_channel       (id_router_053_src_channel),             //          .channel
		.sink_data          (id_router_053_src_data),                //          .data
		.sink_startofpacket (id_router_053_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_053_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_053_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_053_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_053_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_053_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_053_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_053_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_053_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_053_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_053_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_053_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_053_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_053_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_053_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_053_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_053_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_053_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_053_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_053_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_053_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_053_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_053_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_053_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_053_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_053_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_002 rsp_xbar_demux_054 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_008_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_054_src_ready),               //      sink.ready
		.sink_channel       (id_router_054_src_channel),             //          .channel
		.sink_data          (id_router_054_src_data),                //          .data
		.sink_startofpacket (id_router_054_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_054_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_054_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_054_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_054_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_054_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_054_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_054_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_054_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_054_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_054_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_054_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_054_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_054_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_054_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_054_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_054_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_054_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_054_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_054_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_054_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_054_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_054_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_054_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_054_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_054_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_054_src3_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_055 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_055_src_ready),               //      sink.ready
		.sink_channel       (id_router_055_src_channel),             //          .channel
		.sink_data          (id_router_055_src_data),                //          .data
		.sink_startofpacket (id_router_055_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_055_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_055_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_055_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_055_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_055_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_055_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_055_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_055_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_056 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_056_src_ready),               //      sink.ready
		.sink_channel       (id_router_056_src_channel),             //          .channel
		.sink_data          (id_router_056_src_data),                //          .data
		.sink_startofpacket (id_router_056_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_056_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_056_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_056_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_056_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_056_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_056_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_056_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_056_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux rsp_xbar_demux_057 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_057_src_ready),               //      sink.ready
		.sink_channel       (id_router_057_src_channel),             //          .channel
		.sink_data          (id_router_057_src_data),                //          .data
		.sink_startofpacket (id_router_057_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_057_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_057_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_057_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_057_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_057_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_057_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_057_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_057_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_057_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_057_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_057_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_057_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_057_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_057_src1_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_058 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_058_src_ready),               //      sink.ready
		.sink_channel       (id_router_058_src_channel),             //          .channel
		.sink_data          (id_router_058_src_data),                //          .data
		.sink_startofpacket (id_router_058_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_058_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_058_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_058_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_058_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_058_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_058_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_058_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_058_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_059 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_059_src_ready),               //      sink.ready
		.sink_channel       (id_router_059_src_channel),             //          .channel
		.sink_data          (id_router_059_src_data),                //          .data
		.sink_startofpacket (id_router_059_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_059_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_059_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_059_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_059_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_059_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_059_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_059_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_059_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_060 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_060_src_ready),               //      sink.ready
		.sink_channel       (id_router_060_src_channel),             //          .channel
		.sink_data          (id_router_060_src_data),                //          .data
		.sink_startofpacket (id_router_060_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_060_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_060_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_060_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_060_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_060_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_060_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_060_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_060_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_061 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_061_src_ready),               //      sink.ready
		.sink_channel       (id_router_061_src_channel),             //          .channel
		.sink_data          (id_router_061_src_data),                //          .data
		.sink_startofpacket (id_router_061_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_061_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_061_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_061_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_061_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_061_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_061_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_061_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_061_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_062 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_062_src_ready),               //      sink.ready
		.sink_channel       (id_router_062_src_channel),             //          .channel
		.sink_data          (id_router_062_src_data),                //          .data
		.sink_startofpacket (id_router_062_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_062_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_062_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_062_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_062_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_062_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_062_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_062_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_062_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_063 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_063_src_ready),               //      sink.ready
		.sink_channel       (id_router_063_src_channel),             //          .channel
		.sink_data          (id_router_063_src_data),                //          .data
		.sink_startofpacket (id_router_063_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_063_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_063_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_063_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_063_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_063_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_063_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_063_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_063_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_064 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_064_src_ready),               //      sink.ready
		.sink_channel       (id_router_064_src_channel),             //          .channel
		.sink_data          (id_router_064_src_data),                //          .data
		.sink_startofpacket (id_router_064_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_064_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_064_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_064_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_064_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_064_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_064_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_064_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_064_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_demux_001 rsp_xbar_demux_065 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_065_src_ready),               //      sink.ready
		.sink_channel       (id_router_065_src_channel),             //          .channel
		.sink_data          (id_router_065_src_data),                //          .data
		.sink_startofpacket (id_router_065_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_065_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_065_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_065_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_065_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_065_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_065_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_065_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_065_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux rsp_xbar_mux (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid            (rsp_xbar_mux_src_valid),                //          .valid
		.src_data             (rsp_xbar_mux_src_data),                 //          .data
		.src_channel          (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket    (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_017_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_017_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_017_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_017_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_017_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_017_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_018_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_018_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_018_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_018_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_018_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_018_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_019_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_019_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_019_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_019_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_019_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_019_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_020_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_021_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_022_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_023_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_024_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_017_src2_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_017_src2_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_017_src2_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_017_src2_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_017_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_017_src2_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_018_src2_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_018_src2_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_018_src2_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_018_src2_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_018_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_018_src2_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_019_src2_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_019_src2_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_019_src2_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_019_src2_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_019_src2_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_019_src2_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_021_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_021_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_021_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_021_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_021_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_021_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_022_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_022_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_022_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_022_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_022_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_022_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_023_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_023_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_023_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_023_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_023_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_023_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_024_src1_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_024_src1_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_024_src1_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_024_src1_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_024_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_024_src1_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_025_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_025_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_026_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_026_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_027_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_027_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_028_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_002 rsp_xbar_mux_003 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_014_src1_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_014_src1_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_014_src1_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_014_src1_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_014_src1_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_015_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_015_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_015_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_015_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_015_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_016_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_016_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_016_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_016_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_016_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_016_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_022_src2_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_022_src2_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_022_src2_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_022_src2_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_022_src2_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_022_src2_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_023_src2_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_023_src2_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_023_src2_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_023_src2_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_023_src2_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_023_src2_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_024_src2_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_024_src2_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_024_src2_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_024_src2_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_024_src2_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_024_src2_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_029_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_029_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_029_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_030_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_030_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_030_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_030_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_031_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_031_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_031_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_031_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_031_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_032_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_032_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_032_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_032_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_032_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_033_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_033_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_004 rsp_xbar_mux_004 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_004_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_004_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_004_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_014_src2_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_014_src2_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_014_src2_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_014_src2_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_014_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_014_src2_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_015_src2_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_015_src2_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_015_src2_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_015_src2_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_015_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_015_src2_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_016_src2_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_016_src2_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_016_src2_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_016_src2_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_016_src2_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_016_src2_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_022_src3_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_022_src3_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_022_src3_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_022_src3_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_022_src3_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_022_src3_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_023_src3_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_023_src3_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_023_src3_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_023_src3_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_023_src3_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_023_src3_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_024_src3_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_024_src3_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_024_src3_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_024_src3_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_024_src3_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_024_src3_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_030_src1_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_030_src1_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_030_src1_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_030_src1_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_030_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_030_src1_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_031_src1_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_031_src1_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_031_src1_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_031_src1_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_031_src1_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_031_src1_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_032_src1_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_032_src1_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_032_src1_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_032_src1_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_032_src1_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_032_src1_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_033_src1_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_033_src1_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_033_src1_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_033_src1_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_033_src1_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_033_src1_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_034_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_034_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_035_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_035_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_036_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_036_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_037_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_037_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_002 rsp_xbar_mux_005 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_005_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_005_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_005_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_011_src1_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_011_src1_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_011_src1_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_011_src1_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_011_src1_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_012_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_012_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_012_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_012_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_012_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_013_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_013_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_013_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_013_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_013_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_031_src2_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_031_src2_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_031_src2_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_031_src2_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_031_src2_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_031_src2_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_032_src2_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_032_src2_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_032_src2_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_032_src2_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_032_src2_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_032_src2_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_033_src2_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_033_src2_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_033_src2_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_033_src2_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_033_src2_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_033_src2_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_038_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_038_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_038_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_038_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_038_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_039_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_039_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_039_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_039_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_039_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_040_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_040_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_040_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_040_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_040_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_041_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_041_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_041_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_041_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_041_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_042_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_042_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_004 rsp_xbar_mux_006 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_006_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_006_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_006_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_011_src2_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_011_src2_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_011_src2_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_011_src2_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_011_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_011_src2_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_012_src2_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_012_src2_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_012_src2_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_012_src2_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_012_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_012_src2_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_013_src2_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_013_src2_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_013_src2_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_013_src2_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_013_src2_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_013_src2_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_031_src3_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_031_src3_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_031_src3_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_031_src3_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_031_src3_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_031_src3_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_032_src3_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_032_src3_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_032_src3_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_032_src3_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_032_src3_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_032_src3_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_033_src3_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_033_src3_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_033_src3_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_033_src3_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_033_src3_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_033_src3_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_039_src1_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_039_src1_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_039_src1_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_039_src1_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_039_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_039_src1_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_040_src1_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_040_src1_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_040_src1_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_040_src1_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_040_src1_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_040_src1_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_041_src1_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_041_src1_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_041_src1_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_041_src1_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_041_src1_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_041_src1_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_042_src1_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_042_src1_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_042_src1_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_042_src1_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_042_src1_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_042_src1_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_043_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_043_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_044_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_044_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_045_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_045_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_046_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_046_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_002 rsp_xbar_mux_007 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_007_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_007_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_007_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_040_src2_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_040_src2_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_040_src2_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_040_src2_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_040_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_040_src2_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_041_src2_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_041_src2_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_041_src2_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_041_src2_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_041_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_041_src2_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_042_src2_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_042_src2_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_042_src2_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_042_src2_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_042_src2_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_042_src2_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_047_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_047_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_047_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_047_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_047_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_048_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_048_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_048_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_048_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_048_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_049_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_049_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_049_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_049_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_049_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_050_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_050_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_050_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_050_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_050_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_051_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_051_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_051_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_051_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_051_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_052_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_052_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_052_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_052_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_052_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_053_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_053_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_053_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_053_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_053_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_054_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_054_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_054_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_054_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_054_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_054_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_001 rsp_xbar_mux_008 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_008_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_008_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_040_src3_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_040_src3_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_040_src3_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_040_src3_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_040_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_040_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_041_src3_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_041_src3_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_041_src3_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_041_src3_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_041_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_041_src3_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_042_src3_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_042_src3_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_042_src3_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_042_src3_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_042_src3_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_042_src3_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_048_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_048_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_048_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_048_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_048_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_048_src1_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_052_src1_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_052_src1_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_052_src1_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_052_src1_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_052_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_052_src1_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_053_src1_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_053_src1_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_053_src1_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_053_src1_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_053_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_053_src1_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_054_src1_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_054_src1_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_054_src1_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_054_src1_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_054_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_054_src1_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_055_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_055_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_055_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_055_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_055_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_055_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_004 rsp_xbar_mux_009 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_009_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_009_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_009_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_002_src1_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_003_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_004_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_005_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_005_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_006_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_006_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_007_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_007_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_007_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_007_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_008_src1_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_008_src1_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_009_src1_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_009_src1_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_010_src1_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_010_src1_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_010_src1_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_010_src1_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_052_src2_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_052_src2_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_052_src2_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_052_src2_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_052_src2_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_052_src2_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_053_src2_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_053_src2_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_053_src2_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_053_src2_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_053_src2_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_053_src2_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_054_src2_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_054_src2_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_054_src2_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_054_src2_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_054_src2_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_054_src2_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_056_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_056_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_056_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_056_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_056_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_056_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_057_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_057_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_057_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_057_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_057_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_057_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_010 rsp_xbar_mux_010 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_010_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_010_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_010_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_010_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_010_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_010_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_002_src2_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_002_src2_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_002_src2_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_002_src2_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_003_src2_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_003_src2_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_003_src2_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_003_src2_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_003_src2_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_004_src2_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_004_src2_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_004_src2_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_004_src2_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_004_src2_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_004_src2_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_005_src2_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_005_src2_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_005_src2_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_005_src2_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_005_src2_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_005_src2_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_006_src2_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_006_src2_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_006_src2_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_006_src2_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_006_src2_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_006_src2_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_007_src2_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_007_src2_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_007_src2_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_007_src2_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_007_src2_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_007_src2_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_008_src2_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_008_src2_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_008_src2_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_008_src2_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_008_src2_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_008_src2_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_009_src2_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_009_src2_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_009_src2_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_009_src2_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_009_src2_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_009_src2_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_010_src2_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_010_src2_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_010_src2_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_010_src2_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_010_src2_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_052_src3_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_052_src3_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_052_src3_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_052_src3_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_052_src3_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_052_src3_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_053_src3_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_053_src3_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_053_src3_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_053_src3_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_053_src3_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_053_src3_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_054_src3_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_054_src3_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_054_src3_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_054_src3_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_054_src3_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_054_src3_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_057_src1_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_057_src1_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_057_src1_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_057_src1_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_057_src1_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_057_src1_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_058_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_058_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_058_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_058_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_058_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_058_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_059_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_059_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_059_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_059_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_059_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_059_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_060_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_060_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_060_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_060_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_060_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_060_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_061_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_061_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_061_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_061_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_061_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_061_src0_endofpacket)    //          .endofpacket
	);

	SoC_rsp_xbar_mux_011 rsp_xbar_mux_011 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_011_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_011_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_011_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_011_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_011_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_011_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_002_src3_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_002_src3_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_002_src3_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_002_src3_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_003_src3_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_003_src3_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_003_src3_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_003_src3_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_003_src3_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_004_src3_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_004_src3_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_004_src3_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_004_src3_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_004_src3_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_004_src3_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_005_src3_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_005_src3_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_005_src3_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_005_src3_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_005_src3_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_005_src3_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_006_src3_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_006_src3_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_006_src3_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_006_src3_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_006_src3_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_006_src3_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_007_src3_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_007_src3_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_007_src3_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_007_src3_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_007_src3_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_007_src3_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_008_src3_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_008_src3_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_008_src3_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_008_src3_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_008_src3_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_008_src3_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_009_src3_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_009_src3_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_009_src3_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_009_src3_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_009_src3_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_009_src3_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_010_src3_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_010_src3_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_010_src3_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_010_src3_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_010_src3_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_010_src3_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_011_src3_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_011_src3_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_011_src3_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_011_src3_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_011_src3_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_011_src3_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_012_src3_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_012_src3_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_012_src3_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_012_src3_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_012_src3_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_012_src3_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_013_src3_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_013_src3_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_013_src3_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_013_src3_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_013_src3_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_013_src3_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_014_src3_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_014_src3_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_014_src3_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_014_src3_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_014_src3_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_014_src3_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_015_src3_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_015_src3_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_015_src3_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_015_src3_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_015_src3_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_015_src3_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_016_src3_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_016_src3_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_016_src3_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_016_src3_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_016_src3_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_016_src3_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_017_src3_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_017_src3_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_017_src3_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_017_src3_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_017_src3_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_017_src3_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_018_src3_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_018_src3_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_018_src3_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_018_src3_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_018_src3_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_018_src3_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_019_src3_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_019_src3_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_019_src3_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_019_src3_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_019_src3_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_019_src3_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_062_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_062_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_062_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_062_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_062_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_062_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_063_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_063_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_063_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_063_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_063_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_063_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_064_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_064_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_064_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_064_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_064_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_064_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_065_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_065_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_065_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_065_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_065_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_065_src0_endofpacket)    //          .endofpacket
	);

	SoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),       // receiver8.irq
		.sender_irq    (cpu_0_d_irq_irq)                 //    sender.irq
	);

	SoC_irq_mapper_001 irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_001_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_001_receiver6_irq),       // receiver6.irq
		.sender_irq    (cpu_1_d_irq_irq)                     //    sender.irq
	);

	SoC_irq_mapper_002 irq_mapper_002 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_002_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_002_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_001_receiver6_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_002_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu_2_d_irq_irq)                     //    sender.irq
	);

	SoC_irq_mapper_003 irq_mapper_003 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_004_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_003_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_003_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_003_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_002_receiver4_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_003_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver6_irq),           // receiver5.irq
		.sender_irq    (cpu_3_d_irq_irq)                     //    sender.irq
	);

	SoC_irq_mapper_003 irq_mapper_004 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_005_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_004_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_004_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_004_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_003_receiver4_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_004_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver7_irq),           // receiver5.irq
		.sender_irq    (cpu_4_d_irq_irq)                     //    sender.irq
	);

	SoC_irq_mapper_005 irq_mapper_005 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_006_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_005_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_005_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_005_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_004_receiver4_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver8_irq),           // receiver4.irq
		.sender_irq    (cpu_5_d_irq_irq)                     //    sender.irq
	);

endmodule
